// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. 
// LAST TIME SAVED: Nov 20 19:10:52 2014
// NETLIST TIME: Nov 21 11:04:30 2014

module aibcr3_esd ( io );

inout  io;



endmodule


