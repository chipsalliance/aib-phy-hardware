// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. All rights reserved
// ==========================================================================
//
// Module name    : aib_ioring
// Description    : Behavioral model of AIB io buffers
// Revision       : 1.0
// ============================================================================
module aib_ioring 
 #(
    parameter DATAWIDTH = 20
    )
(
inout wire  [DATAWIDTH-1:0]     iopad_txdat, 
inout wire  [DATAWIDTH-1:0]     iopad_rxdat, 
inout wire             iopad_txclkb, 
inout wire             iopad_txclk,
inout wire             iopad_txfck, 
inout wire             iopad_txfckb,
inout wire             iopad_stck, 
inout wire             iopad_stckb,
inout wire             iopad_stl, 
inout wire             iopad_std,
inout wire             iopad_rstno, 
inout wire             iopad_arstno,
inout wire             iopad_spareo, 
inout wire             iopad_sparee,
inout wire             iopad_rxclkb, 
inout wire             iopad_rxclk,
inout wire             iopad_rxfckb, 
inout wire             iopad_rxfck,
inout wire             iopad_srckb, 
inout wire             iopad_srck,
inout wire             iopad_srl, 
inout wire             iopad_srd,
inout wire             iopad_rstni, 
inout wire             iopad_arstni,

input          tx_launch_clk, //Clock for SDR/DDR data, output data clock,ns_fwd_clk_frmac
output wire    fs_rvc_clk_tomac, //rxclki originally
output wire    fs_fwd_clk_tomac, //rxfcki originally
input          ns_rvc_clk_frmac, //txfcko originally
input          dig_rstb, //reset for io buffer
input          iddren,
input          idataselb, //output async data selection
input          itxen,
input [2:0]    irxen,
input [DATAWIDTH-1:0]   idat0,
input [DATAWIDTH-1:0]   idat1,
output wire [DATAWIDTH-1:0]     data_out0,
output wire [DATAWIDTH-1:0]     data_out1,
input       std_out,
input       stl_out,
output wire srd_in,
output wire srl_in,
output wire sr_clk_in,
input       sr_clk_out,
input       adapter_rstno,
input       rstn_out,
output wire adapter_rstni,
output wire rstn_in,

input                  jtag_clkdr_in, 
output wire            scan_out,
input                  jtag_intest,
input                  jtag_mode_in,
input                  jtag_rstb, //reset for io buffer
input                  jtag_rstb_en,
input                  jtag_weakpdn,
input                  jtag_weakpu,
input                  jtag_tx_scanen_in,
input                  scan_in,

input       [DATAWIDTH-1:0]     tx_shift_en,
input       [DATAWIDTH-1:0]     rx_shift_en,
input                  shift_en_txclkb,
input                  shift_en_txfckb,
input                  shift_en_stckb,
input                  shift_en_stl,
input                  shift_en_arstno,
input                  shift_en_txclk,
input                  shift_en_std,
input                  shift_en_stck,
input                  shift_en_txfck,
input                  shift_en_rstno,
input                  shift_en_rxclkb,
input                  shift_en_rxfckb,
input                  shift_en_srckb,
input                  shift_en_srl,
input                  shift_en_arstni,
input                  shift_en_rxclk,
input                  shift_en_rxfck,
input                  shift_en_srck,
input                  shift_en_srd,
input                  shift_en_rstni,

input       idataselb_arstno,
input       idataselb_rstno,
input       idataselb_stck,
input       idataselb_std,
input       idataselb_stl,

input     vccl_aib,
input     vssl_aib );


wire         idat0_std, idat1_std;
wire         idat0_stl, idat1_stl;
wire         pcs_data_out0_rxfck;
wire         odat_async_srd;
wire         odat_async_srl;
wire         odat_async_srck;
wire         idat0_stck, idat0_stckb;
wire         rx_distclk;
wire         rx_strbclk;

wire  [DATAWIDTH-1:0]     idat0_poutp; 
wire  [DATAWIDTH-1:0]     idat1_poutp; 

wire  [2:0] irxen_spareo;
wire        itxen_spareo;
wire        odat_async_spareo;

wire  [2:0] irxen_sparee;
wire        itxen_sparee;
wire        odat_async_sparee;

wire        rxfcki;
wire        rxclki;

wire        rxclk_rstb, rxclkb_rstb;

wire        txfcko;

assign      txfcko = iddren ? tx_launch_clk : ~tx_launch_clk;

assign rxclk_rstb = shift_en_rxclk ? dig_rstb  : vccl_aib;
assign rxclkb_rstb = shift_en_rxclkb ? dig_rstb  : vccl_aib;

assign fs_fwd_clk_tomac = rxfcki;

assign fs_rvc_clk_tomac = rxclki;
assign idat0_std = std_out;
assign idat1_std = idat0_std;

assign idat0_stl = stl_out;
assign idat1_stl = idat0_stl;

assign srd_in = odat_async_srd;
assign srl_in = odat_async_srl;

assign sr_clk_in = odat_async_srck;
assign idat0_stck = sr_clk_out;
assign idat0_stckb = ~sr_clk_out;

//assign rx_distclk = rxclki;
//assign rx_strbclk = rxclki;

assign rx_distclk = rxfcki;
assign rx_strbclk = rxfcki;

assign irxen_spareo[2:0] = shift_en_arstno ? {vssl_aib, vccl_aib,vssl_aib} : irxen[2:0];
assign itxen_spareo = shift_en_arstno ?  vccl_aib : vssl_aib;

assign irxen_sparee[2:0] = shift_en_rstno ? {vssl_aib, vccl_aib,vssl_aib} : irxen[2:0];
assign itxen_sparee = shift_en_rstno ?  vccl_aib : vssl_aib;

wire [DATAWIDTH-1:0] nc_oclk, nc_oclkb, nc_odat0;
wire [DATAWIDTH-1:0] nc_odat_async, nc_odat_async_aib_pout, nc_odat1_aib_pout, nc_oclk_aib_pout;
wire [DATAWIDTH-1:0] nc_oclkn_pout, nc_oclkb_aib_pout, nc_odat0_aib_pout, nc_odat1;
wire [DATAWIDTH-1:0] nc_async_dat_pinpi, nc_idat1_pinp, nc_idat0_pinp, nc_oclk_pinp;
wire [DATAWIDTH-1:0] jtag_clkdr_outn_pinp, nc_oclkb_pinp, nc_odat_async_pinp;
wire [DATAWIDTH-1:0] pcs_data_out0_pinp, pcs_data_out1_pinp;

wire [DATAWIDTH-1:0] nc_async_dat_poutp, jtag_clkdr_outn_poutp;
wire [DATAWIDTH-1:0] nc_async_dat_pinp, nc_odat_async_out0_pinp, nc_oclkb_out0_pinp;
wire [DATAWIDTH-1:0] nc_oclk_out0_pinp, nc_oclkn_out0_pinp;

wire [DATAWIDTH-1:0] jtag_rx_scan_out_rxdat;
wire [DATAWIDTH:0] jtag_rx_scan_out_poutp;

assign jtag_rx_scan_out_poutp[DATAWIDTH]= jtag_tx_scanen_in;

if (DATAWIDTH >20) 
begin
aib_buffx1_top txdat19 ( .idata1_in1_jtag_out(idat1_poutp[19]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp19),
     .idata0_in1_jtag_out(idat0_poutp[19]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp19),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .dig_rstb(dig_rstb),
     .oclk_out(nc_oclk[19]), .oclkb_out(nc_oclkb[19]),
     .odat0_out(nc_odat0[19]), .odat1_out(nc_odat1[19]),
     .odat_async_out(nc_odat_async[19]), 
     .async_dat_in0(vssl_aib), .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp19),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[19]),
     .idata0_in1(idat0_poutp[21]), .idata1_in0(idat1[19]),
     .idata1_in1(idat1_poutp[21]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp19), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[19]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[19]), 
     .odat1_aib(nc_odat1_aib_pout[19]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[19]),
     .odat0_aib(nc_odat0_aib_pout[19]),
     .oclk_aib(nc_oclk_aib_pout[19]),
     .oclkb_aib(nc_oclkb_aib_pout[19]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[20]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[19]), .oclkn(nc_oclkn_pout[19]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
end
else
begin
aib_buffx1_top txdat19 ( .idata1_in1_jtag_out(idat1_poutp[19]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp19),
     .idata0_in1_jtag_out(idat0_poutp[19]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp19),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .dig_rstb(dig_rstb),
     .oclk_out(nc_oclk[19]), .oclkb_out(nc_oclkb[19]),
     .odat0_out(nc_odat0[19]), .odat1_out(nc_odat1[19]),
     .odat_async_out(nc_odat_async[19]), 
     .async_dat_in0(vssl_aib), .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp19),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[19]),
     .idata0_in1(vssl_aib), .idata1_in0(idat1[19]),
     .idata1_in1(vssl_aib), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp19), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[19]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[19]), 
     .odat1_aib(nc_odat1_aib_pout[19]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[19]),
     .odat0_aib(nc_odat0_aib_pout[19]),
     .oclk_aib(nc_oclk_aib_pout[19]),
     .oclkb_aib(nc_oclkb_aib_pout[19]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[20]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[19]), .oclkn(nc_oclkn_pout[19]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
end


aib_buffx1_top txdat17 ( .idata1_in1_jtag_out(idat1_poutp[17]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp17),
     .idata0_in1_jtag_out(idat0_poutp[17]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp17),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[17]),
     .oclkb_out(nc_oclkb[17]), .odat0_out(nc_odat0[17]),
     .odat1_out(nc_odat1[17]), .odat_async_out(nc_odat_async[17]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp17),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[17]),
     .idata0_in1(idat0_poutp[19]), .idata1_in0(idat1[17]),
     .idata1_in1(idat1_poutp[19]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp17), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[17]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[17]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[17]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[17]),
     .odat0_aib(nc_odat0_aib_pout[17]),
     .oclk_aib(nc_oclk_aib_pout[17]),
     .oclkb_aib(nc_oclkb_aib_pout[17]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[18]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[17]), .oclkn(nc_oclkn_pout[17]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txdat15 ( .idata1_in1_jtag_out(idat1_poutp[15]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp15),
     .idata0_in1_jtag_out(idat0_poutp[15]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp15),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[15]),
     .oclkb_out(nc_oclkb[15]), .odat0_out(nc_odat0[15]),
     .odat1_out(nc_odat1[15]), .odat_async_out(nc_odat_async[15]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp15),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[15]),
     .idata0_in1(idat0_poutp[17]), .idata1_in0(idat1[15]),
     .idata1_in1(idat1_poutp[17]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp15), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[15]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[15]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[15]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[15]),
     .odat0_aib(nc_odat0_aib_pout[15]),
     .oclk_aib(nc_oclk_aib_pout[15]),
     .oclkb_aib(nc_oclkb_aib_pout[15]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[16]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[15]), .oclkn(nc_oclkn_pout[15]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txdat13 ( .idata1_in1_jtag_out(idat1_poutp[13]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp13),
     .idata0_in1_jtag_out(idat0_poutp[13]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp13),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[13]),
     .oclkb_out(nc_oclkb[13]), .odat0_out(nc_odat0[13]),
     .odat1_out(nc_odat1[13]), .odat_async_out(nc_odat_async[13]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp13),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[13]),
     .idata0_in1(idat0_poutp[15]), .idata1_in0(idat1[13]),
     .idata1_in1(idat1_poutp[15]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp13), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[13]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[13]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[13]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[13]),
     .odat0_aib(nc_odat0_aib_pout[13]),
     .oclk_aib(nc_oclk_aib_pout[13]),
     .oclkb_aib(nc_oclkb_aib_pout[13]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[14]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[13]), .oclkn(nc_oclkn_pout[13]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));


aib_buffx1_top txdat11 ( .idata1_in1_jtag_out(idat1_poutp[11]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp11),
     .idata0_in1_jtag_out(idat0_poutp[11]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp11),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[11]),
     .oclkb_out(nc_oclkb[11]), .odat0_out(nc_odat0[11]),
     .odat1_out(nc_odat1[11]), .odat_async_out(nc_odat_async[11]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp11),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[11]),
     .idata0_in1(idat0_poutp[13]), .idata1_in0(idat1[11]),
     .idata1_in1(idat1_poutp[13]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp11), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[11]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[11]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[11]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[11]),
     .odat0_aib(nc_odat0_aib_pout[11]),
     .oclk_aib(nc_oclk_aib_pout[11]),
     .oclkb_aib(nc_oclkb_aib_pout[11]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[12]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[11]), .oclkn(nc_oclkn_pout[11]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txclkb ( .idata1_in1_jtag_out(idata1_in1_txclkb),
     .async_dat_in1_jtag_out(nc_async_dat_txclkb),
     .idata0_in1_jtag_out(idata0_in1_txclkb),
     .jtag_clkdr_outn(jtag_clkdr_outn_txclkb),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk_txclkb),
     .oclkb_out(nc_oclkb_txclkb), .odat0_out(nc_odat0_txclkb),
     .odat1_out(nc_odat1_txclkb), .odat_async_out(nc_odat_async_txclkb),
     .async_dat_in0(~ns_rvc_clk_frmac),
     .async_dat_in1(~ns_rvc_clk_frmac),
     .iclkin_dist_in0(jtag_clkdr_outn_txclkb),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(~ns_rvc_clk_frmac),
     //.idata0_in1(idat0_poutp[11]), .idata1_in0(~ns_rvc_clk_frmac),
     //.idata1_in1(idat1_poutp[11]), .idataselb_in0(vccl_aib),
     .idata0_in1(idat0_poutp[1]), .idata1_in0(~ns_rvc_clk_frmac),
     .idata1_in1(idat1_poutp[1]), .idataselb_in0(vccl_aib),
     .idataselb_in1(idataselb), .iddren_in0(vccl_aib),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_txclkb), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_txclkb),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(shift_en_txclkb), 
     //.dig_rstb(dig_rstb),
     .dig_rstb(vccl_aib),
     .odat1_aib(nc_odat1_aib_txclkb),
     .jtag_rx_scan_out(jtag_rx_scan_out_txclkb),
     .odat0_aib(nc_odat0_aib_txclkb),
     .oclk_aib(nc_oclk_aib_txclkb),
     .oclkb_aib(nc_oclkb_aib_txclkb), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     //.jtag_tx_scan_in(jtag_rx_scan_out_poutp[10]),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[0]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txclkb), .oclkn(nc_oclkn_txclkb),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txdat9 ( .idata1_in1_jtag_out(idat1_poutp[9]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp9),
     .idata0_in1_jtag_out(idat0_poutp[9]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp9),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[9]),
     .oclkb_out(nc_oclkb[9]), .odat0_out(nc_odat0[9]),
     .odat1_out(nc_odat1[9]), .odat_async_out(nc_odat_async[9]),
     .async_dat_in0(~txfcko),
     .async_dat_in1(~txfcko),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp9),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[9]),
     .idata0_in1(idata0_in1_txclkb), .idata1_in0(idat1[9]),
     .idata1_in1(idata1_in1_txclkb), .idataselb_in0(idataselb),
     .idataselb_in1(vccl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp9), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[9]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[9]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[9]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[9]),
     .odat0_aib(nc_odat0_aib_pout[9]), .oclk_aib(nc_oclk_aib_pout[9]),
     .oclkb_aib(nc_oclkb_aib_pout[9]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_txclk),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[9]), .oclkn(nc_oclkn_pout[9]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txdat7 ( .idata1_in1_jtag_out(idat1_poutp[7]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp7),
     .idata0_in1_jtag_out(idat0_poutp[7]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp7),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[7]),
     .oclkb_out(nc_oclkb[7]), .odat0_out(nc_odat0[7]),
     .odat1_out(nc_odat1[7]), .odat_async_out(nc_odat_async[7]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp7),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[7]),
     .idata0_in1(idat0_poutp[9]), .idata1_in0(idat1[7]),
     .idata1_in1(idat1_poutp[9]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp7), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[7]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[7]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[7]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[7]),
     .odat0_aib(nc_odat0_aib_pout[7]), .oclk_aib(nc_oclk_aib_pout[7]),
     .oclkb_aib(nc_oclkb_aib_pout[7]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[8]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[7]), .oclkn(nc_oclkn_pout[7]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txdat5 ( .idata1_in1_jtag_out(idat1_poutp[5]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp5),
     .idata0_in1_jtag_out(idat0_poutp[5]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp5),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[5]),
     .oclkb_out(nc_oclkb[5]), .odat0_out(nc_odat0[5]),
     .odat1_out(nc_odat1[5]), .odat_async_out(nc_odat_async[5]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp5),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[5]),
     .idata0_in1(idat0_poutp[7]), .idata1_in0(idat1[5]),
     .idata1_in1(idat1_poutp[7]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp5), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[5]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[5]), 
     .dig_rstb(dig_rstb), 
     .odat1_aib(nc_odat1_aib_pout[5]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[5]),
     .odat0_aib(nc_odat0_aib_pout[5]), .oclk_aib(nc_oclk_aib_pout[5]),
     .oclkb_aib(nc_oclkb_aib_pout[5]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[6]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[5]), .oclkn(nc_oclkn_pout[5]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txdat3 ( .idata1_in1_jtag_out(idat1_poutp[3]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp3),
     .idata0_in1_jtag_out(idat0_poutp[3]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp3),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[3]),
     .oclkb_out(nc_oclkb[3]), .odat0_out(nc_odat0[3]),
     .odat1_out(nc_odat1[3]), .odat_async_out(nc_odat_async[3]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp3),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[3]),
     .idata0_in1(idat0_poutp[5]), .idata1_in0(idat1[3]),
     .idata1_in1(idat1_poutp[5]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp3), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[3]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[3]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[3]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[3]),
     .odat0_aib(nc_odat0_aib_pout[3]), .oclk_aib(nc_oclk_aib_pout[3]),
     .oclkb_aib(nc_oclkb_aib_pout[3]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[4]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[3]), .oclkn(nc_oclkn_pout[3]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txdat1 ( .idata1_in1_jtag_out(idat1_poutp[1]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp1),
     .idata0_in1_jtag_out(idat0_poutp[1]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp1),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk[1]), .oclkb_out(nc_oclkb[1]),
     .odat0_out(nc_odat0[1]), .odat1_out(nc_odat1[1]),
     .odat_async_out(nc_odat_async[1]), 
     .async_dat_in0(vssl_aib), .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp1),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[1]),
     .idata0_in1(idat0_poutp[3]), .idata1_in0(idat1[1]),
     .idata1_in1(idat1_poutp[3]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp1), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[1]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[1]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[1]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[1]),
     .odat0_aib(nc_odat0_aib_pout[1]), .oclk_aib(nc_oclk_aib_pout[1]),
     .oclkb_aib(nc_oclkb_aib_pout[1]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[2]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[1]), .oclkn(nc_oclkn_pout[1]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txfckb ( .idata1_in1_jtag_out(idata1_in1_txfckb),
     .async_dat_in1_jtag_out(nc_async_dat_txfckb),
     .idata0_in1_jtag_out(idata0_in1_txfckb),
     .jtag_clkdr_outn(jtag_clkdr_outn_txfckb),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk_txfckb),
     .oclkb_out(nc_oclkb_txfckb), .odat0_out(nc_odat0_txfckb),
     .odat1_out(nc_odat1_txfckb), .odat_async_out(nc_odat_async_txfckb),
     //.async_dat_in0(~tx_launch_clk),
     //.async_dat_in1(~tx_launch_clk),
     .async_dat_in0(~txfcko),
     .async_dat_in1(~txfcko),
     .iclkin_dist_in0(jtag_clkdr_outn_txfckb),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(~tx_launch_clk),
     //.idata0_in1(idat0_poutp[1]), .idata1_in0(~tx_launch_clk),
     //.idata1_in1(idat1_poutp[1]), .idataselb_in0(vccl_aib),
     .idata0_in1(idat0_poutp[11]), .idata1_in0(~tx_launch_clk),
     .idata1_in1(idat1_poutp[11]), .idataselb_in0(vccl_aib),
     .idataselb_in1(idataselb), .iddren_in0(vccl_aib),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_txfckb), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_txfckb),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(shift_en_txfckb), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_txfckb),
     .jtag_rx_scan_out(jtag_rx_scan_out_txfckb),
     .odat0_aib(nc_odat0_aib_txfckb),
     .oclk_aib(nc_oclk_aib_txfckb),
     .oclkb_aib(nc_oclkb_aib_txfckb), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     //.jtag_tx_scan_in(jtag_rx_scan_out_poutp[0]),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[10]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txfckb), .oclkn(nc_oclkn_txfckb),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top stckb ( .idata1_in1_jtag_out(idata1_in1_stckb),
     .async_dat_in1_jtag_out(nc_async_dat_stckb),
     .idata0_in1_jtag_out(idata0_in1_stckb),
     .jtag_clkdr_outn(jtag_clkdr_outn_stckb),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk_stckb),
     .oclkb_out(nc_oclkb_stckb), .odat0_out(nc_odat0_stckb),
     .odat1_out(nc_odat1_stckb), .odat_async_out(nc_odat_async_stckb),
     .async_dat_in0(idat0_stckb),
     .async_dat_in1(idata0_in1_txclkb),
     .iclkin_dist_in0(jtag_clkdr_outn_stckb),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0_stckb),
     .idata0_in1(idata0_in1_txclkb), .idata1_in0(idat0_stckb),
     .idata1_in1(idata1_in1_txclkb), .idataselb_in0(idataselb_stck),
     .idataselb_in1(vccl_aib), .iddren_in0(vccl_aib),
     .iddren_in1(vccl_aib), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_stckb), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_stckb),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(shift_en_stckb), 
     //.dig_rstb(dig_rstb),
     .dig_rstb(vccl_aib),
     .odat1_aib(nc_odat1_aib_stckb),
     .jtag_rx_scan_out(jtag_rx_scan_out_stckb),
     .odat0_aib(nc_odat0_aib_stckb),
     .oclk_aib(nc_oclk_aib_stckb),
     .oclkb_aib(nc_oclkb_aib_stckb), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_txfck),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_stckb), .oclkn(nc_oclkn_stckb),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top stl ( .idata1_in1_jtag_out(idata1_in1_stl),
     .async_dat_in1_jtag_out(nc_async_dat_stl),
     .idata0_in1_jtag_out(idata0_in1_stl),
     .jtag_clkdr_outn(jtag_clkdr_outn_stl),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk_stl),
     .oclkb_out(nc_oclkb_stl), .odat0_out(nc_odat0_stl),
     .odat1_out(nc_odat1_stl), .odat_async_out(nc_odat_async_stl),
     .async_dat_in0(idat0_stl),
     .async_dat_in1(idata0_in1_stckb),
     .iclkin_dist_in0(jtag_clkdr_outn_stl),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0_stl),
     .idata0_in1(idata0_in1_stckb), .idata1_in0(idat1_stl),
     .idata1_in1(idata1_in1_stckb), .idataselb_in0(idataselb_stl),
     .idataselb_in1(vccl_aib), .iddren_in0(vccl_aib),
     .iddren_in1(vccl_aib), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_stl), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_stl),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(shift_en_stl), 
     //.dig_rstb(dig_rstb),
     .dig_rstb(vccl_aib),
     .odat1_aib(nc_odat1_aib_stl),
     .jtag_rx_scan_out(jtag_rx_scan_out_stl),
     .odat0_aib(nc_odat0_aib_stl),
     .oclk_aib(nc_oclk_aib_stl),
     .oclkb_aib(nc_oclkb_aib_stl), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_stck),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_stl), .oclkn(nc_oclkn_stl),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top arstno ( .idata1_in1_jtag_out(idata1_in1_arstno),
     .async_dat_in1_jtag_out(nc_async_dat_arstno),
     .idata0_in1_jtag_out(idata0_in1_arstno),
     .jtag_clkdr_outn(jtag_clkdr_outn_arstno),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk_arstno),
     .oclkb_out(nc_oclkb_arstno), .odat0_out(nc_odat0_arstno),
     .odat1_out(nc_odat1_arstno), .odat_async_out(nc_odat_async_arstno),
     .async_dat_in0(adapter_rstno),
     .async_dat_in1(idata0_in1_stl),
     .iclkin_dist_in0(jtag_clkdr_outn_arstno),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(adapter_rstno),
     .idata0_in1(idata0_in1_stl), .idata1_in0(vccl_aib),
     .idata1_in1(idata1_in1_stl), .idataselb_in0(idataselb_arstno),
     .idataselb_in1(vccl_aib), .iddren_in0(vccl_aib),
     .iddren_in1(vccl_aib), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_arstno), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_arstno),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(shift_en_arstno), 
     //.dig_rstb(dig_rstb),
     .dig_rstb(vccl_aib),
     .odat1_aib(nc_odat1_aib_arstno),
     .jtag_rx_scan_out(jtag_rx_scan_out_arstno),
     .odat0_aib(nc_odat0_aib_arstno),
     .oclk_aib(nc_oclk_aib_arstno),
     .oclkb_aib(nc_oclkb_aib_arstno), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_std),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_arstno), .oclkn(nc_oclkn_arstno),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top spareo ( .idata1_in1_jtag_out(idata1_in1_spareo),
     .async_dat_in1_jtag_out(nc_async_dat_spareo),
     .idata0_in1_jtag_out(idata0_in1_spareo),
     .jtag_clkdr_outn(jtag_clkdr_outn_spareo),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk_spareo),
     .oclkb_out(nc_oclkb_spareo), .odat0_out(nc_odat0_spareo),
     .odat1_out(nc_odat1_spareo), .odat_async_out(odat_async_spareo),
     .async_dat_in0(adapter_rstno),
     .async_dat_in1(adapter_rstno),
     .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk), .idata0_in0(adapter_rstno),
     .idata0_in1(adapter_rstno), .idata1_in0(adapter_rstno),
     .idata1_in1(adapter_rstno), .idataselb_in0(idataselb_arstno),
     .idataselb_in1(idataselb_arstno), .iddren_in0(vccl_aib),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0(irxen_spareo[2:0]),
     .irxen_in1(irxen_spareo[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(itxen_spareo), .itxen_in1(itxen_spareo), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_spareo),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(vssl_aib), 
     //.dig_rstb(dig_rstb),
     .dig_rstb(vccl_aib),
     .odat1_aib(odat1_aib_spareo),
     .jtag_rx_scan_out(jtag_rx_scan_out_spareo),
     .odat0_aib(odat0_aib_spareo),
     .oclk_aib(nc_oclk_aib_spareo),
     .oclkb_aib(nc_oclkb_aib_spareo), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_rstno),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_spareo), .oclkn(nc_oclkn_spareo),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));


if (DATAWIDTH >20) 
begin
aib_buffx1_top txdat18 ( .idata1_in1_jtag_out(idat1_poutp[18]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp18),
     .idata0_in1_jtag_out(idat0_poutp[18]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp18),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[18]),
     .oclkb_out(nc_oclkb[18]), .odat0_out(nc_odat0[18]),
     .odat1_out(nc_odat1[18]), .odat_async_out(nc_odat_async[18]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp18),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[18]),
     .idata0_in1(idat0_poutp[20]), .idata1_in0(idat1[18]),
     .idata1_in1(idat1_poutp[20]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp18), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[18]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[18]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[18]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[18]),
     .odat0_aib(nc_odat0_aib_pout[18]),
     .oclk_aib(nc_oclk_aib_pout[18]),
     .oclkb_aib(nc_oclkb_aib_pout[18]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[19]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[18]), .oclkn(nc_oclkn_pout[18]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
end
else 
begin
aib_buffx1_top txdat18 ( .idata1_in1_jtag_out(idat1_poutp[18]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp18),
     .idata0_in1_jtag_out(idat0_poutp[18]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp18),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[18]),
     .oclkb_out(nc_oclkb[18]), .odat0_out(nc_odat0[18]),
     .odat1_out(nc_odat1[18]), .odat_async_out(nc_odat_async[18]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp18),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[18]),
     .idata0_in1(vssl_aib), .idata1_in0(idat1[18]),
     .idata1_in1(vssl_aib), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp18), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[18]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[18]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[18]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[18]),
     .odat0_aib(nc_odat0_aib_pout[18]),
     .oclk_aib(nc_oclk_aib_pout[18]),
     .oclkb_aib(nc_oclkb_aib_pout[18]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[19]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[18]), .oclkn(nc_oclkn_pout[18]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
end

aib_buffx1_top txdat16 ( .idata1_in1_jtag_out(idat1_poutp[16]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp16),
     .idata0_in1_jtag_out(idat0_poutp[16]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp16),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[16]),
     .oclkb_out(nc_oclkb[16]), .odat0_out(nc_odat0[16]),
     .odat1_out(nc_odat1[16]), .odat_async_out(nc_odat_async[16]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp16),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[16]),
     .idata0_in1(idat0_poutp[18]), .idata1_in0(idat1[16]),
     .idata1_in1(idat1_poutp[18]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp16), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[16]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[16]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[16]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[16]),
     .odat0_aib(nc_odat0_aib_pout[16]),
     .oclk_aib(nc_oclk_aib_pout[16]),
     .oclkb_aib(nc_oclkb_aib_pout[16]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[17]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[16]), .oclkn(nc_oclkn_pout[16]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txdat14 ( .idata1_in1_jtag_out(idat1_poutp[14]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp14),
     .idata0_in1_jtag_out(idat0_poutp[14]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp14),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[14]),
     .oclkb_out(nc_oclkb[14]), .odat0_out(nc_odat0[14]),
     .odat1_out(nc_odat1[14]), .odat_async_out(nc_odat_async[14]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp14),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[14]),
     .idata0_in1(idat0_poutp[16]), .idata1_in0(idat1[14]),
     .idata1_in1(idat1_poutp[16]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp14), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[14]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[14]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[14]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[14]),
     .odat0_aib(nc_odat0_aib_pout[14]),
     .oclk_aib(nc_oclk_aib_pout[14]),
     .oclkb_aib(nc_oclkb_aib_pout[14]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[15]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[14]), .oclkn(nc_oclkn_pout[14]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txdat12 ( .idata1_in1_jtag_out(idat1_poutp[12]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp12),
     .idata0_in1_jtag_out(idat0_poutp[12]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp12),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[12]),
     .oclkb_out(nc_oclkb[12]), .odat0_out(nc_odat0[12]),
     .odat1_out(nc_odat1[12]), .odat_async_out(nc_odat_async[12]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp12),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[12]),
     .idata0_in1(idat0_poutp[14]), .idata1_in0(idat1[12]),
     .idata1_in1(idat1_poutp[14]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp12), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[12]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[12]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[12]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[12]),
     .odat0_aib(nc_odat0_aib_pout[12]),
     .oclk_aib(nc_oclk_aib_pout[12]),
     .oclkb_aib(nc_oclkb_aib_pout[12]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[13]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[12]), .oclkn(nc_oclkn_pout[12]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txdat10 ( .idata1_in1_jtag_out(idat1_poutp[10]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp10),
     .idata0_in1_jtag_out(idat0_poutp[10]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp10),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[10]),
     .oclkb_out(nc_oclkb[10]), .odat0_out(nc_odat0[10]),
     .odat1_out(nc_odat1[10]), .odat_async_out(nc_odat_async[10]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp10),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[10]),
     .idata0_in1(idat0_poutp[12]), .idata1_in0(idat1[10]),
     .idata1_in1(idat1_poutp[12]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp10), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[10]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[10]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[10]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[10]),
     .odat0_aib(nc_odat0_aib_pout[10]),
     .oclk_aib(nc_oclk_aib_pout[10]),
     .oclkb_aib(nc_oclkb_aib_pout[10]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[11]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[10]), .oclkn(nc_oclkn_pout[10]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txclk ( .idata1_in1_jtag_out(idata1_in1_txclk),
     .async_dat_in1_jtag_out(nc_async_dat_txclk),
     .idata0_in1_jtag_out(idata0_in1_txclk),
     .jtag_clkdr_outn(jtag_clkdr_outn_txclk),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk_txclk),
     .oclkb_out(nc_oclkb_txclk), .odat0_out(nc_odat0_txclk),
     .odat1_out(nc_odat1_txclk), .odat_async_out(nc_odat_async_txclk),
     .async_dat_in0(ns_rvc_clk_frmac),
     .async_dat_in1(ns_rvc_clk_frmac),
     .iclkin_dist_in0(jtag_clkdr_outn_txclk),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(ns_rvc_clk_frmac),
     //.idata0_in1(idat0_poutp[10]), .idata1_in0(ns_rvc_clk_frmac),
     //.idata1_in1(idat1_poutp[10]), .idataselb_in0(vccl_aib),
     .idata0_in1(idat0_poutp[0]), .idata1_in0(ns_rvc_clk_frmac),
     .idata1_in1(idat1_poutp[0]), .idataselb_in0(vccl_aib),
     .idataselb_in1(idataselb), .iddren_in0(vccl_aib),
     .iddren_in1(iddren), .ilaunch_clk_in0(ns_rvc_clk_frmac),
     .ilaunch_clk_in1(ns_rvc_clk_frmac), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_txclk), .istrbclk_in1(vssl_aib),
     .itxen_in0(vccl_aib), .itxen_in1(vccl_aib), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_txclk),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(shift_en_txclk), 
     //.dig_rstb(dig_rstb),
     .dig_rstb(vccl_aib),
     .odat1_aib(nc_odat1_aib_txclk),
     .jtag_rx_scan_out(jtag_rx_scan_out_txclk),
     .odat0_aib(nc_odat0_aib_txclk),
     .oclk_aib(nc_oclk_aib_txclk),
     .oclkb_aib(nc_oclkb_aib_txclk), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_txclkb),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txclk), .oclkn(nc_oclkn_txclk),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txdat8 ( .idata1_in1_jtag_out(idat1_poutp[8]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp8),
     .idata0_in1_jtag_out(idat0_poutp[8]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp8),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[8]),
     .oclkb_out(nc_oclkb[8]), .odat0_out(nc_odat0[8]),
     .odat1_out(nc_odat1[8]), .odat_async_out(nc_odat_async[8]),
     .async_dat_in0(txfcko),
     .async_dat_in1(txfcko),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp8),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[8]),
     .idata0_in1(idata0_in1_txfck), .idata1_in0(idat1[8]),
     .idata1_in1(idata1_in1_txfck), .idataselb_in0(idataselb),
     .idataselb_in1(vccl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp8), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[8]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[8]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[8]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[8]),
     .odat0_aib(nc_odat0_aib_pout[8]), .oclk_aib(nc_oclk_aib_pout[8]),
     .oclkb_aib(nc_oclkb_aib_pout[8]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[9]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[8]), .oclkn(nc_oclkn_pout[8]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txdat6 ( .idata1_in1_jtag_out(idat1_poutp[6]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp6),
     .idata0_in1_jtag_out(idat0_poutp[6]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp6),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[6]),
     .oclkb_out(nc_oclkb[6]), .odat0_out(nc_odat0[6]),
     .odat1_out(nc_odat1[6]), .odat_async_out(nc_odat_async[6]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp6),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[6]),
     .idata0_in1(idat0_poutp[8]), .idata1_in0(idat1[6]),
     .idata1_in1(idat1_poutp[8]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp6), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[6]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[6]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[6]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[6]),
     .odat0_aib(nc_odat0_aib_pout[6]), .oclk_aib(nc_oclk_aib_pout[6]),
     .oclkb_aib(nc_oclkb_aib_pout[6]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[7]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[6]), .oclkn(nc_oclkn_pout[6]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txdat4 ( .idata1_in1_jtag_out(idat1_poutp[4]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp4),
     .idata0_in1_jtag_out(idat0_poutp[4]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp4),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[4]),
     .oclkb_out(nc_oclkb[4]), .odat0_out(nc_odat0[4]),
     .odat1_out(nc_odat1[4]), .odat_async_out(nc_odat_async[4]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp4),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[4]),
     .idata0_in1(idat0_poutp[6]), .idata1_in0(idat1[4]),
     .idata1_in1(idat1_poutp[6]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp4), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[4]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[4]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[4]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[4]),
     .odat0_aib(nc_odat0_aib_pout[4]), .oclk_aib(nc_oclk_aib_pout[4]),
     .oclkb_aib(nc_oclkb_aib_pout[4]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[5]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[4]), .oclkn(nc_oclkn_pout[4]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txdat2 ( .idata1_in1_jtag_out(idat1_poutp[2]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp2),
     .idata0_in1_jtag_out(idat0_poutp[2]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp2),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[2]),
     .oclkb_out(nc_oclkb[2]), .odat0_out(nc_odat0[2]),
     .odat1_out(nc_odat1[2]), .odat_async_out(nc_odat_async[2]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp2),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[2]),
     .idata0_in1(idat0_poutp[4]), .idata1_in0(idat1[2]),
     .idata1_in1(idat1_poutp[4]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp2), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[2]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[2]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[2]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[2]),
     .odat0_aib(nc_odat0_aib_pout[2]), .oclk_aib(nc_oclk_aib_pout[2]),
     .oclkb_aib(nc_oclkb_aib_pout[2]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[3]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[2]), .oclkn(nc_oclkn_pout[2]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txdat0 ( .idata1_in1_jtag_out(idat1_poutp[0]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp0),
     .idata0_in1_jtag_out(idat0_poutp[0]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp0),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk[0]), .oclkb_out(nc_oclkb[0]),
     .odat0_out(nc_odat0[0]), .odat1_out(nc_odat1[0]),
     .odat_async_out(nc_odat_async[0]), 
     .async_dat_in0(vssl_aib), .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp0),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[0]),
     .idata0_in1(idat0_poutp[2]), .idata1_in0(idat1[0]),
     .idata1_in1(idat1_poutp[2]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib,
     vccl_aib, vssl_aib}), .irxen_in1({vssl_aib,vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_poutp0), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen),
     .oclk_in1(vssl_aib), .odat_async_aib(odat_async_pout0),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[0]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[0]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[0]),
     .odat0_aib(nc_odat0_aib_pout[0]), .oclk_aib(nc_oclk_aib_pout[0]),
     .oclkb_aib(nc_oclkb_aib_pout[0]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[1]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[0]), .oclkn(nc_oclkn_pout[0]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top txfck ( .idata1_in1_jtag_out(idata1_in1_txfck),
     .async_dat_in1_jtag_out(nc_async_dat_txfck),
     .idata0_in1_jtag_out(idata0_in1_txfck),
     .jtag_clkdr_outn(jtag_clkdr_outn_txfck),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk_txfck),
     .oclkb_out(nc_oclkb_txfck), .odat0_out(nc_odat0_txfck),
     .odat1_out(nc_odat1_txfck), .odat_async_out(nc_odat_async_txfck),
     //.async_dat_in0(tx_launch_clk),
     //.async_dat_in1(tx_launch_clk),
     .async_dat_in0(txfcko),
     .async_dat_in1(txfcko),
     .iclkin_dist_in0(jtag_clkdr_outn_txfck),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(tx_launch_clk),
     //.idata0_in1(idat0_poutp[0]), .idata1_in0(tx_launch_clk),
     //.idata1_in1(idat1_poutp[0]), .idataselb_in0(vccl_aib),
     .idata0_in1(idat0_poutp[10]), .idata1_in0(tx_launch_clk),
     .idata1_in1(idat1_poutp[10]), .idataselb_in0(vccl_aib),
     .idataselb_in1(idataselb), .iddren_in0(vccl_aib),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_txfck), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_txfck),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(shift_en_txfck), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_txfck),
     .jtag_rx_scan_out(jtag_rx_scan_out_txfck),
     .odat0_aib(nc_odat0_aib_txfck),
     .oclk_aib(nc_oclk_aib_txfck),
     .oclkb_aib(nc_oclkb_aib_txfck), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_txfckb),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txfck), .oclkn(nc_oclkn_txfck),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top stck ( .idata1_in1_jtag_out(idata1_in1_stck),
     .async_dat_in1_jtag_out(nc_async_dat_stck),
     .idata0_in1_jtag_out(idata0_in1_stck),
     .jtag_clkdr_outn(jtag_clkdr_outn_stck),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk_stck),
     .oclkb_out(nc_oclkb_stck), .odat0_out(nc_odat0_stck),
     .odat1_out(nc_odat1_stck), .odat_async_out(nc_odat_async_stck),
     .async_dat_in0(idat0_stck),
     .async_dat_in1(idata0_in1_txclk),
     .iclkin_dist_in0(jtag_clkdr_outn_stck),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0_stck),
     .idata0_in1(idata0_in1_txclk), .idata1_in0(idat0_stck),
     .idata1_in1(idata1_in1_txclk), .idataselb_in0(idataselb_stck),
     .idataselb_in1(vccl_aib), .iddren_in0(vccl_aib),
     .iddren_in1(vccl_aib), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_stck), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_stck),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(shift_en_stck), 
     //.dig_rstb(dig_rstb),
     .dig_rstb(vccl_aib),
     .odat1_aib(nc_odat1_aib_stck),
     .jtag_rx_scan_out(jtag_rx_scan_out_stck),
     .odat0_aib(nc_odat0_aib_stck),
     .oclk_aib(nc_oclk_aib_stck),
     .oclkb_aib(nc_oclkb_aib_stck), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_stckb),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_stck), .oclkn(nc_oclkn_stck),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top std ( .idata1_in1_jtag_out(idata1_in1_std),
     .async_dat_in1_jtag_out(nc_async_dat_std),
     .idata0_in1_jtag_out(idata0_in1_std),
     .jtag_clkdr_outn(jtag_clkdr_outn_std),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk_std),
     .oclkb_out(nc_oclkb_std), .odat0_out(nc_odat0_std),
     .odat1_out(nc_odat1_std), .odat_async_out(nc_odat_async_std),
     .async_dat_in0(idat0_std),
     .async_dat_in1(idata0_in1_stck),
     .iclkin_dist_in0(jtag_clkdr_outn_std),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0_std),
     .idata0_in1(idata0_in1_stck), .idata1_in0(idat1_std),
     .idata1_in1(idata1_in1_stck), .idataselb_in0(idataselb_std),
     .idataselb_in1(vccl_aib), .iddren_in0(vccl_aib),
     .iddren_in1(vccl_aib), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_std), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_std),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(shift_en_std), 
     //.dig_rstb(dig_rstb),
     .dig_rstb(vccl_aib),
     .odat1_aib(nc_odat1_aib_std),
     .jtag_rx_scan_out(jtag_rx_scan_out_std),
     .odat0_aib(nc_odat0_aib_std),
     .oclk_aib(nc_oclk_aib_std),
     .oclkb_aib(nc_oclkb_aib_std), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_stl),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_std), .oclkn(nc_oclkn_std),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top rstno ( .idata1_in1_jtag_out(idata1_in1_rstno),
     .async_dat_in1_jtag_out(nc_async_dat_rstno),
     .idata0_in1_jtag_out(idata0_in1_rstno),
     .jtag_clkdr_outn(jtag_clkdr_outn_rstno),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk_rstno),
     .oclkb_out(nc_oclkb_rstno), .odat0_out(nc_odat0_rstno),
     .odat1_out(nc_odat1_rstno), .odat_async_out(nc_odat_async_rstno),
     .async_dat_in0(rstn_out),
     .async_dat_in1(idata0_in1_std),
     .iclkin_dist_in0(jtag_clkdr_outn_rstno),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(rstn_out),
     .idata0_in1(idata0_in1_std), .idata1_in0(vccl_aib),
     .idata1_in1(idata1_in1_std), .idataselb_in0(idataselb_rstno),
     .idataselb_in1(vccl_aib), .iddren_in0(vccl_aib),
     .iddren_in1(vccl_aib), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(jtag_clkdr_outn_rstno), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_rstno),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(shift_en_rstno), 
     //.dig_rstb(dig_rstb),
     .dig_rstb(vccl_aib),
     .odat1_aib(nc_odat1_aib_rstno),
     .jtag_rx_scan_out(jtag_rx_scan_out_rstno),
     .odat0_aib(nc_odat0_aib_rstno),
     .oclk_aib(nc_oclk_aib_rstno),
     .oclkb_aib(nc_oclkb_aib_rstno), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_arstno),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_rstno), .oclkn(nc_oclkn_rstno),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top sparee ( .idata1_in1_jtag_out(idata1_in1_sparee),
     .async_dat_in1_jtag_out(nc_async_dat_sparee),
     .idata0_in1_jtag_out(idata0_in1_sparee),
     .jtag_clkdr_outn(jtag_clkdr_outn_sparee),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk_sparee),
     .oclkb_out(nc_oclkb_sparee), .odat0_out(nc_odat0_sparee),
     .odat1_out(nc_odat1_sparee), .odat_async_out(odat_async_sparee),
     .async_dat_in0(rstn_out),
     .async_dat_in1(rstn_out),
     .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk), .idata0_in0(rstn_out),
     .idata0_in1(rstn_out), .idata1_in0(rstn_out),
     .idata1_in1(rstn_out), .idataselb_in0(idataselb_rstno),
     .idataselb_in1(idataselb_rstno), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0(irxen_sparee[2:0]),
     .irxen_in1(irxen_sparee[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(itxen_sparee), .itxen_in1(itxen_sparee), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_sparee),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(vssl_aib), 
     //.dig_rstb(dig_rstb),
     .dig_rstb(vccl_aib),
     .odat1_aib(odat1_aib_sparee),
     .jtag_rx_scan_out(jtag_rx_scan_out_sparee),
     .odat0_aib(odat0_aib_sparee),
     .oclk_aib(nc_oclk_aib_sparee),
     .oclkb_aib(nc_oclkb_aib_sparee), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_spareo),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_sparee), .oclkn(nc_oclkn_sparee),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));


aib_buffx1_top rxdat19 ( .idata1_in1_jtag_out(nc_idat1_pinp19),
     .async_dat_in1_jtag_out(nc_async_dat_pinp19),
     .idata0_in1_jtag_out(nc_idat0_pinp19),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp19),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp19), .oclkb_out(nc_oclkb_pinp19),
     .odat0_out(data_out0[19]),
     .odat1_out(data_out1[19]),
     .odat_async_out(nc_odat_async_pinp19),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib), .idata0_in1(vssl_aib),
     .idata1_in0(vssl_aib), .idata1_in1(vssl_aib),
     .idataselb_in0(vccl_aib), .idataselb_in1(vssl_aib),
     .iddren_in0(iddren), .iddren_in1(iddren),
     .ilaunch_clk_in0(vssl_aib), .ilaunch_clk_in1(vssl_aib),
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk),
     .istrbclk_in1(rx_strbclk), .itxen_in0(vssl_aib),
     .itxen_in1(vssl_aib), .oclk_in1(vssl_aib),
     .odat_async_aib(odirectin_data_pinp19), .oclkb_in1(vssl_aib),
     .odat0_in1(pcs_data_out0_pinp17),
     .odat1_in1(pcs_data_out1_pinp17), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[19]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(pcs_data_out1_pinp[19]),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[19]),
     .odat0_aib(pcs_data_out0_pinp[19]), .oclk_aib(ncdrx_oclk_pinp19),
     .oclkb_aib(ncdrx_oclkb_pinp19),
     .jtag_clkdr_in(jtag_clkdr_in), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[18]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_rxdat[19]), .oclkn(ncdrx_oclkn_pinp19),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxdat17 ( .idata1_in1_jtag_out(nc_idat1_pinp17),
     .async_dat_in1_jtag_out(nc_async_dat_pinp17),
     .idata0_in1_jtag_out(nc_idat0_pinp17),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp17),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp17), .oclkb_out(nc_oclkb_pinp17),
     .odat0_out(data_out0[17]),
     .odat1_out(data_out1[17]),
     .odat_async_out(nc_odat_async_pinp17),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_pinp17),
     .oclkb_in1(vssl_aib), .odat0_in1(ncdrx_odat0_pinp15),
     .odat1_in1(ncdrx_odat1_pinp15), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[17]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(pcs_data_out1_pinp17),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[17]),
     .odat0_aib(pcs_data_out0_pinp17), .oclk_aib(nc_oclk_out0_pinp17),
     .oclkb_aib(nc_oclkb_out0_pinp17), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[16]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxdat[17]),
     .oclkn(nc_oclkn_out0_pinp17), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxdat15 ( .idata1_in1_jtag_out(nc_idat1_pinp15),
     .async_dat_in1_jtag_out(nc_async_dat_pinp15),
     .idata0_in1_jtag_out(nc_idat0_pinp15),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp15),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp15), .oclkb_out(nc_oclkb_pinp15),
     .odat0_out(data_out0[15]),
     .odat1_out(data_out1[15]),
     .odat_async_out(nc_odat_async_pinp15),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_pinp15),
     .oclkb_in1(vssl_aib), .odat0_in1(pcs_data_out0_pinp13),
     .odat1_in1(pcs_data_out1_pinp13), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[15]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(ncdrx_odat1_pinp15),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[15]),
     .odat0_aib(ncdrx_odat0_pinp15), .oclk_aib(ncdrx_oclk_pinp15),
     .oclkb_aib(ncdrx_oclkb_pinp15),
     .jtag_clkdr_in(jtag_clkdr_in), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[14]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxdat[15]),
     .oclkn(ncdrx_oclkn_pinp15), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxdat13 ( .idata1_in1_jtag_out(nc_idat1_pinp13),
     .async_dat_in1_jtag_out(nc_async_dat_pinp13),
     .idata0_in1_jtag_out(nc_idat0_pinp13),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp13),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp13), .oclkb_out(nc_oclkb_pinp13),
     .odat0_out(data_out0[13]),
     .odat1_out(data_out1[13]),
     .odat_async_out(nc_odat_async_pinp13),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_pinp13),
     .oclkb_in1(vssl_aib), .odat0_in1(pcs_data_out0_pinp11),
     .odat1_in1(pcs_data_out1_pinp11), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[13]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(pcs_data_out1_pinp13),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[13]),
     .odat0_aib(pcs_data_out0_pinp13), .oclk_aib(nc_oclk_out0_pinp13),
     .oclkb_aib(nc_oclkb_out0_pinp13), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[12]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxdat[13]),
     .oclkn(nc_oclkn_out0_pinp13), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxdat11 ( .idata1_in1_jtag_out(nc_idat1_pinp11),
     .async_dat_in1_jtag_out(nc_async_dat_pinp11),
     .idata0_in1_jtag_out(nc_idat0_pinp11),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp11),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp11), .oclkb_out(nc_oclkb_pinp11),
     .odat0_out(data_out0[11]),
     .odat1_out(data_out1[11]),
     .odat_async_out(nc_odat_async_pinp11),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_pinp11),
     .oclkb_in1(vssl_aib), .odat0_in1(pcs_data_out0_rxfckb),
     .odat1_in1(pcs_data_out1_rxfckb), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[11]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(pcs_data_out1_pinp11),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[11]),
     .odat0_aib(pcs_data_out0_pinp11), .oclk_aib(nc_oclk_out0_pinp11),
     .oclkb_aib(nc_oclkb_out0_pinp11), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[10]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxdat[11]),
     .oclkn(nc_oclkn_out0_pinp11), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxclkb ( .idata1_in1_jtag_out(nc_idat1_rxclkb),
     .async_dat_in1_jtag_out(nc_async_dat_rxclkb),
     .idata0_in1_jtag_out(nc_idat0_rxclkb),
     .jtag_clkdr_outn(jtag_clkdr_outn_rxclkb),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_rxclkb), .oclkb_out(nc_oclkb_rxclkb),
     .odat0_out(data_out0_rxclkb),
     .odat1_out(data_out1_rxclkb),
     .odat_async_out(nc_odat_async_rxclkb),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vccl_aib), .iddren_in0(vccl_aib),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_rxclkb),
     //.oclkb_in1(vssl_aib), .odat0_in1(ncdrx_odat0_pinp9),
     //.odat1_in1(ncdrx_odat1_pinp9), .odat_async_in1(vssl_aib),
     .oclkb_in1(vssl_aib), .odat0_in1(pcs_data_out0_srckb),
     .odat1_in1(pcs_data_out1_srckb), .odat_async_in1(nc_odat_async_out0_srckb),
     .shift_en(shift_en_rxclkb), 
     //.dig_rstb(dig_rstb),
     //.dig_rstb(vccl_aib),
     .dig_rstb(rxclkb_rstb),
     .odat1_aib(pcs_data_out1_rxclkb),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxclkb),
     .odat0_aib(pcs_data_out0_rxclkb), .oclk_aib(nc_oclk_out0_rxclkb),
     .oclkb_aib(nc_oclkb_out0_rxclkb), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_rxclk),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxclkb),
     .oclkn(nc_oclkn_out0_rxclkb), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxdat9 ( .idata1_in1_jtag_out(nc_idat1_pinp9),
     .async_dat_in1_jtag_out(nc_async_dat_pinp9),
     .idata0_in1_jtag_out(nc_idat0_pinp9),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp9),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp9), .oclkb_out(nc_oclkb_pinp9),
     .odat0_out(data_out0[9]), .odat1_out(data_out1[9]),
     .odat_async_out(nc_odat_async_pinp9),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vccl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk),
     .istrbclk_in1(vssl_aib), .itxen_in0(vssl_aib),
     .itxen_in1(vssl_aib), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_out0_pinp9), .oclkb_in1(vssl_aib),
     .odat0_in1(pcs_data_out0_pinp7), .odat1_in1(pcs_data_out1_pinp7),
     .odat_async_in1(vssl_aib), .shift_en(rx_shift_en[9]),
     .dig_rstb(dig_rstb),
     .odat1_aib(ncdrx_odat1_pinp9),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[9]),
     .odat0_aib(ncdrx_odat0_pinp9), .oclk_aib(ncdrx_oclk_pinp9),
     .oclkb_aib(ncdrx_oclkb_pinp9),
     .jtag_clkdr_in(jtag_clkdr_in), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[8]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxdat[9]),
     .oclkn(oclkn_pinp9), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxdat7 ( .idata1_in1_jtag_out(nc_idat1_pinp7),
     .async_dat_in1_jtag_out(nc_async_dat_pinp7),
     .idata0_in1_jtag_out(nc_idat0_pinp7),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp7),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp7), .oclkb_out(nc_oclkb_pinp7),
     .odat0_out(data_out0[7]), .odat1_out(data_out1[7]),
     .odat_async_out(nc_odat_async_pinp7),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_pinp7),
     .oclkb_in1(vssl_aib), .odat0_in1(ncdrx_odat0_pinp5),
     .odat1_in1(ncdrx_odat1_pinp5), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[7]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(pcs_data_out1_pinp7),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[7]),
     .odat0_aib(pcs_data_out0_pinp7), .oclk_aib(nc_oclk_out0_pinp7),
     .oclkb_aib(nc_oclkb_out0_pinp7),
     .jtag_clkdr_in(jtag_clkdr_in), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[6]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxdat[7]),
     .oclkn(nc_oclkn_out0_pinp7), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxdat5 ( .idata1_in1_jtag_out(nc_idat1_pinp5),
     .async_dat_in1_jtag_out(nc_async_dat_pinp5),
     .idata0_in1_jtag_out(nc_idat0_pinp5),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp5),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp5), .oclkb_out(nc_oclkb_pinp5),
     .odat0_out(data_out0[5]), .odat1_out(data_out1[5]),
     .odat_async_out(nc_odat_async_pinp5),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_pinp5),
     .oclkb_in1(vssl_aib), .odat0_in1(pcs_data_out0_pinp3),
     .odat1_in1(pcs_data_out1_pinp3), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[5]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(ncdrx_odat1_pinp5),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[5]),
     .odat0_aib(ncdrx_odat0_pinp5), .oclk_aib(ncdrx_oclk_pinp5),
     .oclkb_aib(ncdrx_oclkb_pinp5),
     .jtag_clkdr_in(jtag_clkdr_in), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[4]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .test_weakpd(jtag_weakpdn),
     .test_weakpu(jtag_weakpu), .iopad(iopad_rxdat[5]),
     .oclkn(ncdrx_oclkn_pinp5), .iclkn(vssl_aib));

aib_buffx1_top rxdat3 ( .idata1_in1_jtag_out(nc_idat1_pinp3),
     .async_dat_in1_jtag_out(nc_async_dat_pinp3),
     .idata0_in1_jtag_out(nc_idat0_pinp3),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp3),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp3), .oclkb_out(nc_oclkb_pinp3),
     .odat0_out(data_out0[3]), .odat1_out(data_out1[3]),
     .odat_async_out(nc_odat_async_pinp3),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_pinp3),
     .oclkb_in1(vssl_aib), .odat0_in1(pcs_data_out0_pinp1),
     .odat1_in1(pcs_data_out1_pinp1), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[3]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(pcs_data_out1_pinp3),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[3]),
     .odat0_aib(pcs_data_out0_pinp3), .oclk_aib(nc_oclk_out0_pinp3),
     .oclkb_aib(nc_oclkb_out0_pinp3),
     .jtag_clkdr_in(jtag_clkdr_in), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[2]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxdat[3]),
     .oclkn(nc_oclkn_out0_pinp3), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxdat1 ( .idata1_in1_jtag_out(nc_idat1_pinp1),
     .async_dat_in1_jtag_out(nc_async_dat_pinp1),
     .idata0_in1_jtag_out(nc_idat0_pinp1),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp1),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp1), .oclkb_out(nc_oclkb_pinp1),
     .odat0_out(data_out0[1]), .odat1_out(data_out1[1]),
     .odat_async_out(nc_odat_async_pinp1),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vccl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_pinp1),
     .oclkb_in1(vssl_aib), .odat0_in1(pcs_data_out0_rxclkb),
     .odat1_in1(pcs_data_out1_rxclkb),
     .odat_async_in1(vssl_aib), .shift_en(rx_shift_en[1]),
     .dig_rstb(dig_rstb),
     .odat1_aib(pcs_data_out1_pinp1),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[1]),
     .odat0_aib(pcs_data_out0_pinp1), .oclk_aib(nc_oclk_out0_pinp1),
     .oclkb_aib(nc_oclkb_out0_pinp1),
     .jtag_clkdr_in(jtag_clkdr_in), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[0]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .test_weakpd(jtag_weakpdn),
     .test_weakpu(jtag_weakpu), .iopad(iopad_rxdat[1]),
     .oclkn(nc_oclkn_out0_pinp1), .iclkn(vssl_aib));

aib_buffx1_top rxfckb ( .idata1_in1_jtag_out(nc_idat1_rxfckb),
     .async_dat_in1_jtag_out(nc_async_dat_rxfckb),
     .idata0_in1_jtag_out(nc_idat0_rxfckb),
     .jtag_clkdr_outn(jtag_clkdr_outn_rxfckb),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_rxfckb), .oclkb_out(nc_oclkb_rxfckb),
     .odat0_out(data_out0_rxfckb),
     .odat1_out(data_out1_rxfckb),
     .odat_async_out(nc_odat_async_rxfckb),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(vccl_aib),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_rxfckb),
     //.oclkb_in1(vssl_aib), .odat0_in1(pcs_data_out0_srckb),
     //.odat1_in1(pcs_data_out1_srckb), .odat_async_in1(vssl_aib),
     .oclkb_in1(vssl_aib), .odat0_in1(data_out0[9]),
     .odat1_in1(data_out1[9]), .odat_async_in1(nc_odat_async_out0_pinp9),
     .shift_en(shift_en_rxfckb), 
     .dig_rstb(dig_rstb),
     .odat1_aib(pcs_data_out1_rxfckb),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxfckb),
     .odat0_aib(pcs_data_out0_rxfckb), .oclk_aib(nc_oclk_out0_rxfckb),
     .oclkb_aib(nc_oclkb_out0_rxfckb), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_rxfck),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxfckb),
     .oclkn(nc_oclkn_out0_rxfckb), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top srckb ( .idata1_in1_jtag_out(nc_idat1_srckb),
     .async_dat_in1_jtag_out(nc_async_dat_srckb),
     .idata0_in1_jtag_out(nc_idat0_srckb),
     .jtag_clkdr_outn(jtag_clkdr_outn_srckb),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_srckb), .oclkb_out(nc_oclkb_srckb),
     .odat0_out(pcs_data_out0_srckb),
     .odat1_out(pcs_data_out1_srckb),
     .odat_async_out(nc_odat_async_srckb),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(vccl_aib),
     .iddren_in1(vssl_aib), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_srckb),
     .oclkb_in1(vssl_aib), .odat0_in1(pcs_data_out0_srl),
     .odat1_in1(pcs_data_out1_srckb), .odat_async_in1(nc_odat_async_out0_srl),
     .shift_en(shift_en_srckb), 
     //.dig_rstb(dig_rstb),
     .dig_rstb(vccl_aib),
     .odat1_aib(pcs_data_out1_srckb),
     .jtag_rx_scan_out(jtag_rx_scan_out_srckb),
     .odat0_aib(pcs_data_out0_srckb), .oclk_aib(nc_oclk_out0_srckb),
     .oclkb_aib(nc_oclkb_out0_srckb), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_srck),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_srckb),
     .oclkn(nc_oclkn_out0_srckb), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top srl ( .idata1_in1_jtag_out(nc_idat1_srl),
     .async_dat_in1_jtag_out(nc_async_dat_srl),
     .idata0_in1_jtag_out(nc_idat0_srl),
     .jtag_clkdr_outn(jtag_clkdr_outn_srl),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_srl), .oclkb_out(nc_oclkb_srl),
     .odat0_out(pcs_data_out0_srl),
     .odat1_out(pcs_data_out1_srl),
     .odat_async_out(odat_async_srl),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(vccl_aib),
     .iddren_in1(vssl_aib), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_srl),
     .oclkb_in1(vssl_aib), .odat0_in1(pcs_data_out0_arstni),
     .odat1_in1(pcs_data_out1_arstni), .odat_async_in1(nc_odat_async_out0_arstni),
     .shift_en(shift_en_srl), 
     //.dig_rstb(dig_rstb),
     .dig_rstb(vccl_aib),
     .odat1_aib(pcs_data_out1_srl),
     .jtag_rx_scan_out(jtag_rx_scan_out_srl),
     .odat0_aib(pcs_data_out0_srl), .oclk_aib(nc_oclk_out0_srl),
     .oclkb_aib(nc_oclkb_out0_srl), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_srd),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_srl),
     .oclkn(nc_oclkn_out0_srl), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top arstni ( .idata1_in1_jtag_out(nc_idat1_arstni),
     .async_dat_in1_jtag_out(nc_async_dat_arstni),
     .idata0_in1_jtag_out(nc_idat0_arstni),
     .jtag_clkdr_outn(jtag_clkdr_outn_arstni),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_arstni), .oclkb_out(nc_oclkb_arstni),
     .odat0_out(pcs_data_out0_arstni),
     .odat1_out(pcs_data_out1_arstni),
     .odat_async_out(adapter_rstni),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(vccl_aib),
     .iddren_in1(vssl_aib), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_arstni),
     .oclkb_in1(vssl_aib), .odat0_in1(odat0_aib_sparee),
     .odat1_in1(odat1_aib_sparee), .odat_async_in1(nc_odat_async_aib_sparee),
     .shift_en(shift_en_arstni), 
     //.dig_rstb(dig_rstb),
     .dig_rstb(vccl_aib),
     .odat1_aib(pcs_data_out1_arstni),
     .jtag_rx_scan_out(jtag_rx_scan_out_arstni),
     .odat0_aib(pcs_data_out0_arstni), .oclk_aib(nc_oclk_out0_arstni),
     .oclkb_aib(nc_oclkb_out0_arstni), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_rstni),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_arstni),
     .oclkn(nc_oclkn_out0_arstni), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxdat18 ( .idata1_in1_jtag_out(nc_idat1_pinp18),
     .async_dat_in1_jtag_out(nc_async_dat_pinp18),
     .idata0_in1_jtag_out(nc_idat0_pinp18),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp18),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp18), .oclkb_out(nc_oclkb_pinp18),
     .odat0_out(data_out0[18]),
     .odat1_out(data_out1[18]),
     .odat_async_out(nc_odat_async_pinp18),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib), .idata0_in1(vssl_aib),
     .idata1_in0(vssl_aib), .idata1_in1(vssl_aib),
     .idataselb_in0(vccl_aib), .idataselb_in1(idataselb),
     .iddren_in0(iddren), .iddren_in1(iddren),
     .ilaunch_clk_in0(vssl_aib), .ilaunch_clk_in1(vssl_aib),
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk),
     .istrbclk_in1(vssl_aib), .itxen_in0(vssl_aib),
     .itxen_in1(vssl_aib), .oclk_in1(vssl_aib),
     .odat_async_aib(odirectin_data_pinp18), .oclkb_in1(vssl_aib),
     .odat0_in1(pcs_data_out0_pinp16),
     .odat1_in1(pcs_data_out1_pinp16), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[18]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(pcs_data_out1_pinp[18]),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[18]),
     .odat0_aib(pcs_data_out0_pinp[18]), .oclk_aib(ncdrx_oclk_pinp18),
     .oclkb_aib(ncdrx_oclkb_pinp18),
     .jtag_clkdr_in(jtag_clkdr_in), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[17]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_rxdat[18]), .oclkn(ncdrx_oclkn_pinp18),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxdat16 ( .idata1_in1_jtag_out(nc_idat1_pinp16),
     .async_dat_in1_jtag_out(nc_async_dat_pinp16),
     .idata0_in1_jtag_out(nc_idat0_pinp16),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp16),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp16), .oclkb_out(nc_oclkb_pinp16),
     .odat0_out(data_out0[16]),
     .odat1_out(data_out1[16]),
     .odat_async_out(nc_odat_async_pinp16),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(data_out0[14]),
     .idata0_in1(data_out1[14]), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_pinp16),
     .oclkb_in1(vssl_aib), .odat0_in1(odat0_pinp14),
     .odat1_in1(odat1_pinp14), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[16]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(pcs_data_out1_pinp16),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[16]),
     .odat0_aib(pcs_data_out0_pinp16), .oclk_aib(nc_oclk_out0_pinp16),
     .oclkb_aib(nc_oclkb_out0_pinp16), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[15]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxdat[16]),
     .oclkn(nc_oclkn_out0_pinp16), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxdat14 ( .idata1_in1_jtag_out(nc_idat1_pinp14),
     .async_dat_in1_jtag_out(nc_async_dat_pinp14),
     .idata0_in1_jtag_out(nc_idat0_pinp14),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp14),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp14), .oclkb_out(nc_oclkb_pinp14),
     .odat0_out(data_out0[14]),
     .odat1_out(data_out1[14]),
     .odat_async_out(nc_odat_async_pinp14),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib),
     .odat_async_aib(odirectin_data_out0_pinp14),
     .oclkb_in1(vssl_aib), .odat0_in1(odat0_pinp12),
     .odat1_in1(odat1_pinp12), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[14]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(odat1_pinp14),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[14]),
     .odat0_aib(odat0_pinp14), .oclk_aib(ncdrx_oclk_pinp14),
     .oclkb_aib(ncdrx_oclkb_pinp14),
     .jtag_clkdr_in(jtag_clkdr_in), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[13]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxdat[14]),
     .oclkn(ncdrx_oclkn_pinp14), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxdat12 ( .idata1_in1_jtag_out(nc_idat1_pinp12),
     .async_dat_in1_jtag_out(nc_async_dat_pinp12),
     .idata0_in1_jtag_out(nc_idat0_pinp12),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp12),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp12), .oclkb_out(nc_oclkb_pinp12),
     .odat0_out(data_out0[12]),
     .odat1_out(data_out1[12]),
     .odat_async_out(nc_odat_async_pinp12),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib),
     .odat_async_aib(odirectin_data_out0_pinp12),
     .oclkb_in1(vssl_aib), .odat0_in1(odat0_pinp10),
     .odat1_in1(odat1_pinp10), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[12]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(odat1_pinp12),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[12]),
     .odat0_aib(odat0_pinp12), .oclk_aib(ncdrx_oclkb_out0_pinp12),
     .oclkb_aib(ncdrx_oclkb_out0_pinp12),
     .jtag_clkdr_in(jtag_clkdr_in), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[11]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxdat[12]),
     .oclkn(ncdrx_oclkn_out0_pinp12), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxdat10 ( .idata1_in1_jtag_out(nc_idat1_pinp10),
     .async_dat_in1_jtag_out(nc_async_dat_pinp10),
     .idata0_in1_jtag_out(nc_idat0_pinp10),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp10),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp10), .oclkb_out(nc_oclkb_pinp10),
     .odat0_out(data_out0[10]),
     .odat1_out(data_out1[10]),
     .odat_async_out(nc_odat_async_pinp10),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib),
     .odat_async_aib(odirectin_data_out0_pinp10),
     .oclkb_in1(vssl_aib), .odat0_in1(pcs_data_out0_rxfck),
     .odat1_in1(pcs_data_out1_rxfck), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[10]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(odat1_pinp10),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[10]),
     .odat0_aib(odat0_pinp10), .oclk_aib(ncdrx_oclk_out0_pinp10),
     .oclkb_aib(ncdrx_oclkb_out0_pinp10), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_rxclkb),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxdat[10]),
     .oclkn(ncdrx_oclkn_out0_pinp10), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxclk ( .idata1_in1_jtag_out(nc_idat1_rxclk),
     .async_dat_in1_jtag_out(nc_async_dat_rxclk),
     .idata0_in1_jtag_out(nc_idat0_rxclk),
     .jtag_clkdr_outn(jtag_clkdr_outn_rxclk),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_rxclk), .oclkb_out(nc_oclkb_rxclk),
     .odat0_out(data_out0_rxclk),
     .odat1_out(data_out1_rxclk),
     .odat_async_out(rxclki),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vccl_aib), .iddren_in0(vccl_aib),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(3'b111), .irxen_in1(3'b111),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_rxclk),
     //.oclkb_in1(vssl_aib), .odat0_in1(data_out0[8]),
     //.odat1_in1(data_out1[8]), .odat_async_in1(vssl_aib),
     .oclkb_in1(vssl_aib), .odat0_in1(pcs_data_out0_srck),
     .odat1_in1(pcs_data_out1_srck), .odat_async_in1(nc_odat_async_out0_srck),
     .shift_en(shift_en_rxclk), 
     //.dig_rstb(dig_rstb),
     //.dig_rstb(vccl_aib),
     .dig_rstb(rxclk_rstb),
     .odat1_aib(pcs_data_out1_rxclk),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxclk),
     .odat0_aib(pcs_data_out0_rxclk), .oclk_aib(nc_oclk_out0_rxclk),
     .oclkb_aib(nc_oclkb_out0_rxclk), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     //.jtag_tx_scan_in(jtag_rx_scan_out_rxdat[9]),
     .jtag_tx_scan_in(jtag_rx_scan_out_srckb),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxclk),
     .oclkn(nc_oclkn_out0_rxclk), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxdat8 ( .idata1_in1_jtag_out(nc_idat1_pinp8),
     .async_dat_in1_jtag_out(nc_async_dat_pinp8),
     .idata0_in1_jtag_out(nc_idat0_pinp8),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp8),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp8), .oclkb_out(nc_oclkb_pinp8),
     .odat0_out(data_out0[8]), .odat1_out(data_out1[8]),
     .odat_async_out(nc_odat_async_pinp8),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vccl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_pinp8),
     .oclkb_in1(vssl_aib), .odat0_in1(pcs_data_out0_pinp6),
     .odat1_in1(pcs_data_out1_pinp6), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[8]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(ncdrx_odat1_pinp8),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[8]),
     .odat0_aib(ncdrx_odat0_pinp8), .oclk_aib(oclk_pinp8),
     .oclkb_aib(oclkb_pinp8),
     .jtag_clkdr_in(jtag_clkdr_in), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[7]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxdat[8]),
     .oclkn(ncdrx_oclkn_pinp8), .iclkn(oclkn_pinp9),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxdat6 ( .idata1_in1_jtag_out(nc_idat1_pinp6),
     .async_dat_in1_jtag_out(nc_async_dat_pinp6),
     .idata0_in1_jtag_out(nc_idat0_pinp6),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp6),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp6), .oclkb_out(nc_oclkb_pinp6),
     .odat0_out(data_out0[6]), .odat1_out(data_out1[6]),
     .odat_async_out(nc_odat_async_pinp6),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_pinp6),
     .oclkb_in1(vssl_aib), .odat0_in1(ncdrx_odat0_pinp4),
     .odat1_in1(ncdrx_odat1_pinp4), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[6]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(pcs_data_out1_pinp6),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[6]),
     .odat0_aib(pcs_data_out0_pinp6), .oclk_aib(nc_oclk_out0_pinp6),
     .oclkb_aib(nc_oclkb_out0_pinp6),
     .jtag_clkdr_in(jtag_clkdr_in), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[5]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxdat[6]),
     .oclkn(nc_oclkn_out0_pinp6), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxdat4 ( .idata1_in1_jtag_out(nc_idat1_pinp4),
     .async_dat_in1_jtag_out(nc_async_dat_pinp4),
     .idata0_in1_jtag_out(nc_idat0_pinp4),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp4),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp4), .oclkb_out(nc_oclkb_pinp4),
     .odat0_out(data_out0[4]), .odat1_out(data_out1[4]),
     .odat_async_out(nc_odat_async_pinp4),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_pinp4),
     .oclkb_in1(vssl_aib), .odat0_in1(ncdrx_odat0_out0_pinp2),
     .odat1_in1(ncdrx_odat1_out0_pinp2), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[4]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(ncdrx_odat1_pinp4),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[4]),
     .odat0_aib(ncdrx_odat0_pinp4), .oclk_aib(ncdrx_oclk_pinp4),
     .oclkb_aib(ncdrx_oclkb_pinp4),
     .jtag_clkdr_in(jtag_clkdr_in), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[3]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxdat[4]),
     .oclkn(ncdrx_oclkn_pinp4), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxdat2 ( .idata1_in1_jtag_out(nc_idat1_pinp2),
     .async_dat_in1_jtag_out(nc_async_dat_pinp2),
     .idata0_in1_jtag_out(nc_idat0_pinp2),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp2),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp2), .oclkb_out(nc_oclkb_pinp2),
     .odat0_out(data_out0[2]), .odat1_out(data_out1[2]),
     .odat_async_out(nc_odat_async_pinp2),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(odirectin_data_out0_pinp2),
     .oclkb_in1(vssl_aib), .odat0_in1(ncdrx_odat0_out0_pinp0),
     .odat1_in1(ncdrx_odat1_out0_pinp0), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[2]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(ncdrx_odat1_out0_pinp2),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[2]),
     .odat0_aib(ncdrx_odat0_out0_pinp2),
     .oclk_aib(ncdrx_oclk_out0_pinp2), 
     .oclkb_aib(ncdrx_oclkb_out0_pinp2), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[1]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxdat[2]),
     .oclkn(ncdrx_oclkn_out0_pinp2), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxdat0 ( .idata1_in1_jtag_out(nc_idat1_pinp0),
     .async_dat_in1_jtag_out(nc_async_dat_pinp0),
     .idata0_in1_jtag_out(nc_idat0_pinp0),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp0),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp0), .oclkb_out(nc_oclkb_pinp0),
     .odat0_out(data_out0[0]), .odat1_out(data_out1[0]),
     .odat_async_out(nc_odat_async_pinp0),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(odirectin_data_out0_pinp0),
     .oclkb_in1(vssl_aib), .odat0_in1(pcs_data_out0_rxclk),
     .odat1_in1(pcs_data_out1_rxclk), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[0]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(ncdrx_odat1_out0_pinp0),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[0]),
     .odat0_aib(ncdrx_odat0_out0_pinp0),
     .oclk_aib(ncdrx_oclk_out0_pinp0), 
     .oclkb_aib(ncdrx_oclkb_out0_pinp0), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_rxfckb),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxdat[0]),
     .oclkn(ncdrx_oclkn_out0_pinp0), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rxfck ( .idata1_in1_jtag_out(nc_idat1_rxfck),
     .async_dat_in1_jtag_out(nc_async_dat_rxfck),
     .idata0_in1_jtag_out(nc_idat0_rxfck),
     .jtag_clkdr_outn(jtag_clkdr_outn_rxfck),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_rxfck), .oclkb_out(nc_oclkb_rxfck),
     .odat0_out(data_out0_rxfck),
     .odat1_out(data_out1_rxfck),
     .odat_async_out(rxfcki),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(vccl_aib),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_rxfck),
     .oclkb_in1(vssl_aib), .odat0_in1(data_out0[8]),
     .odat1_in1(data_out1[8]), .odat_async_in1(nc_odat_async_out0_pinp8),
     //.oclkb_in1(vssl_aib), .odat0_in1(pcs_data_out0_srck),
     //.odat1_in1(pcs_data_out1_srck), .odat_async_in1(vssl_aib),
     .shift_en(shift_en_rxfck), 
     .dig_rstb(dig_rstb),
     .odat1_aib(pcs_data_out1_rxfck),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxfck),
     .odat0_aib(pcs_data_out0_rxfck), .oclk_aib(nc_oclk_out0_rxfck),
     .oclkb_aib(nc_oclkb_out0_rxfck), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[9]),
     //.jtag_tx_scan_in(jtag_rx_scan_out_srckb),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxfck),
     .oclkn(nc_oclkn_out0_rxfck), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top srck ( .idata1_in1_jtag_out(nc_idat1_srck),
     .async_dat_in1_jtag_out(nc_async_dat_srck),
     .idata0_in1_jtag_out(nc_idat0_srck),
     .jtag_clkdr_outn(jtag_clkdr_outn_srck),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_srck), .oclkb_out(nc_oclkb_srck),
     .odat0_out(pcs_data_out0_srck),
     .odat1_out(pcs_data_out1_srck),
     .odat_async_out(odat_async_srck),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(vccl_aib),
     .iddren_in1(vssl_aib), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_srck),
     .oclkb_in1(vssl_aib), .odat0_in1(pcs_data_out0_srd),
     .odat1_in1(pcs_data_out1_srd), .odat_async_in1(nc_odat_async_out0_srd),
     .shift_en(shift_en_srck), 
     //.dig_rstb(dig_rstb),
     .dig_rstb(vccl_aib),
     .odat1_aib(pcs_data_out1_srck),
     .jtag_rx_scan_out(jtag_rx_scan_out_srck),
     .odat0_aib(pcs_data_out0_srck), .oclk_aib(nc_oclk_out0_srck),
     .oclkb_aib(nc_oclkb_out0_srck), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_srl),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_srck),
     .oclkn(nc_oclkn_out0_srck), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top srd ( .idata1_in1_jtag_out(nc_idat1_srd),
     .async_dat_in1_jtag_out(nc_async_dat_srd),
     .idata0_in1_jtag_out(nc_idat0_srd),
     .jtag_clkdr_outn(jtag_clkdr_outn_srd),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_srd), .oclkb_out(nc_oclkb_srd),
     .odat0_out(pcs_data_out0_srd),
     .odat1_out(pcs_data_out1_srd),
     .odat_async_out(odat_async_srd),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(vccl_aib),
     .iddren_in1(vssl_aib), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_srd),
     .oclkb_in1(vssl_aib), .odat0_in1(odat0_aib_rstni),
     .odat1_in1(odat1_aib_rstni), .odat_async_in1(nc_odat_async_aib_rstni),
     .shift_en(shift_en_srd), 
     //.dig_rstb(dig_rstb),
     .dig_rstb(vccl_aib),
     .odat1_aib(pcs_data_out1_srd),
     .jtag_rx_scan_out(jtag_rx_scan_out_srd),
     .odat0_aib(pcs_data_out0_srd), .oclk_aib(nc_oclk_out0_srd),
     .oclkb_aib(nc_oclkb_out0_srd), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_arstni),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_srd),
     .oclkn(nc_oclkn_out0_srd), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));

aib_buffx1_top rstni ( .idata1_in1_jtag_out(idata1_in1_rstni),
     .async_dat_in1_jtag_out(nc_async_dat_rstni),
     .idata0_in1_jtag_out(idata0_in1_rstni),
     .jtag_clkdr_outn(jtag_clkdr_outn_rstni),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk_rstni),
     .oclkb_out(nc_oclkb_rstni), .odat0_out(nc_odat0_rstni),
     .odat1_out(nc_odat1_rstni), .odat_async_out(rstn_in),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_rstni),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vccl_aib), .iddren_in0(vssl_aib),
     .iddren_in1(vssl_aib), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0(irxen[2:0]),
     .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_rstni),
     .oclkb_in1(vssl_aib), .odat0_in1(odat0_aib_spareo),
     .odat1_in1(odat1_aib_spareo), .odat_async_in1(nc_odat_async_aib_spareo),
     .shift_en(shift_en_rstni), 
     //.dig_rstb(dig_rstb),
     .dig_rstb(vccl_aib),
     .odat1_aib(odat1_aib_rstni),
     .jtag_rx_scan_out(jtag_rx_scan_out_rstni),
     .odat0_aib(odat0_aib_rstni),
     .oclk_aib(nc_oclk_aib_rstni),
     .oclkb_aib(nc_oclkb_aib_rstni), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_sparee),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_rstni), .oclkn(nc_oclkn_rstni),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));

   genvar i;
   generate
    for (i=20; i<DATAWIDTH; i=i+1) begin:txdatao
     if ((i==DATAWIDTH-1) | (i==DATAWIDTH-2)) begin
aib_buffx1_top txdat ( .idata1_in1_jtag_out(idat1_poutp[i]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp[i]),
     .idata0_in1_jtag_out(idat0_poutp[i]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp[i]),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[i]),
     .oclkb_out(nc_oclkb[i]), .odat0_out(nc_odat0[i]),
     .odat1_out(nc_odat1[i]), .odat_async_out(nc_odat_async[i]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp[i]),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[i]),
     .idata0_in1(vssl_aib), .idata1_in0(idat1[i]),
     .idata1_in1(vssl_aib), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(vssl_aib), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[i]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[i]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[i]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[i]),
     .odat0_aib(nc_odat0_aib_pout[i]),
     .oclk_aib(nc_oclk_aib_pout[i]),
     .oclkb_aib(nc_oclkb_aib_pout[i]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[i+1]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[i]), .oclkn(nc_oclkn_pout[i]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
     end
    else begin
aib_buffx1_top txdat ( .idata1_in1_jtag_out(idat1_poutp[i]),
     .async_dat_in1_jtag_out(nc_async_dat_poutp[i]),
     .idata0_in1_jtag_out(idat0_poutp[i]),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp[i]),
     .jtag_rstb_en(jtag_rstb_en), 
     .jtag_intest(jtag_intest), 
     .oclk_out(nc_oclk[i]),
     .oclkb_out(nc_oclkb[i]), .odat0_out(nc_odat0[i]),
     .odat1_out(nc_odat1[i]), .odat_async_out(nc_odat_async[i]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp[i]),
     .iclkin_dist_in1(vssl_aib), .idata0_in0(idat0[i]),
     .idata0_in1(idat0_poutp[i+2]), .idata1_in0(idat1[i]),
     .idata1_in1(idat1_poutp[i+2]), .idataselb_in0(idataselb),
     .idataselb_in1(idataselb), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk),
     .ilaunch_clk_in1(tx_launch_clk), 
     .irxen_in0({vssl_aib, vccl_aib,
     vssl_aib}), .irxen_in1({vssl_aib, vccl_aib, vssl_aib}),
     .istrbclk_in0(vssl_aib), .istrbclk_in1(vssl_aib),
     .itxen_in0(itxen), .itxen_in1(itxen), .oclk_in1(vssl_aib),
     .odat_async_aib(nc_odat_async_aib_pout[i]),
     .oclkb_in1(vssl_aib), .odat0_in1(vssl_aib),
     .odat1_in1(vssl_aib), .odat_async_in1(vssl_aib),
     .shift_en(tx_shift_en[i]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(nc_odat1_aib_pout[i]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp[i]),
     .odat0_aib(nc_odat0_aib_pout[i]),
     .oclk_aib(nc_oclk_aib_pout[i]),
     .oclkb_aib(nc_oclkb_aib_pout[i]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp[i+1]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), 
     .iopad(iopad_txdat[i]), .oclkn(nc_oclkn_pout[i]),
     .iclkn(vssl_aib), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
    end
    end
   endgenerate



   generate
     for (i=20; i<DATAWIDTH; i=i+1) begin:rxdatai
aib_buffx1_top rxdat ( .idata1_in1_jtag_out(nc_idat1_pinp[i]),
     .async_dat_in1_jtag_out(nc_async_dat_pinp[i]),
     .idata0_in1_jtag_out(nc_idat0_pinp[i]),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp[i]),
     .jtag_rstb_en(jtag_rstb_en),
     .jtag_intest(jtag_intest),
     .oclk_out(nc_oclk_pinp[i]), .oclkb_out(nc_oclkb_pinp[i]),
     .odat0_out(data_out0[i]),
     .odat1_out(data_out1[i]),
     .odat_async_out(nc_odat_async_pinp[i]),
     .async_dat_in0(vssl_aib),
     .async_dat_in1(vssl_aib), .iclkin_dist_in0(rx_distclk),
     .iclkin_dist_in1(rx_distclk),
     .idata0_in0(vssl_aib),
     .idata0_in1(vssl_aib), .idata1_in0(vssl_aib),
     .idata1_in1(vssl_aib), .idataselb_in0(vccl_aib),
     .idataselb_in1(vssl_aib), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(vssl_aib),
     .ilaunch_clk_in1(vssl_aib), 
     .irxen_in0(irxen[2:0]), .irxen_in1(irxen[2:0]),
     .istrbclk_in0(rx_strbclk), .istrbclk_in1(rx_strbclk),
     .itxen_in0(vssl_aib), .itxen_in1(vssl_aib),
     .oclk_in1(vssl_aib), .odat_async_aib(nc_odat_async_out0_pinp[i]),
     .oclkb_in1(vssl_aib), .odat0_in1(pcs_data_out0_pinp[i-2]),
     .odat1_in1(pcs_data_out1_pinp[i-2]), .odat_async_in1(vssl_aib),
     .shift_en(rx_shift_en[i]), 
     .dig_rstb(dig_rstb),
     .odat1_aib(pcs_data_out1_pinp[i]),
     .jtag_rx_scan_out(jtag_rx_scan_out_rxdat[i]),
     .odat0_aib(pcs_data_out0_pinp[i]), .oclk_aib(nc_oclk_out0_pinp[i]),
     .oclkb_aib(nc_oclkb_out0_pinp[i]), .jtag_clkdr_in(jtag_clkdr_in),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_rxdat[i-1]),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .iopad(iopad_rxdat[i]),
     .oclkn(nc_oclkn_out0_pinp[i]), .iclkn(vssl_aib),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
     end
   endgenerate




endmodule

