// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. 
// *****************************************************************************
// *****************************************************************************
// Copyright © 2016 Altera Corporation.                                            
// *****************************************************************************
//  Module Name :  c3lib_dv_defines                                  
//  Date        :  Wed May  4 13:46:15 2016                                 
//  Description :                                                    
// *****************************************************************************

`ifndef __C3LIB_DV_DEFINES__
  `define __C3LIB_DV_DEFINES__

  `define INT_C3LIB_RTL_MODE
  `define FUNCTIONAL


`endif //__C3LIB_DV_DEFINES_V__

