// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. All rights reserved
// ==========================================================================

// This testsbench shows how to connect 24 channel AIB (all channels are independent)
// in loopback mode. DCC/DLL are bypassed. The delay setting is static
// 03/13/2019


`timescale 1ps/1ps

module top;


    //------------------------------------------------------------------------------------------
    // Clock generation
    
    parameter CFG_AVMM_CLK_PERIOD = 4000;
    parameter OSC_CLK_PERIOD      = 1000;
    parameter PMA_CLK_PERIOD      = 1000;
        
    reg   i_cfg_avmm_clk = 1'b0;
    reg	  i_osc_clk = 1'b0;
    reg   i_rx_pma_clk = 1'b0;
    reg   i_rx_pma_div2_clk = 1'b0;
    reg   i_tx_pma_clk = 1'b0;
       
      //clock gen
      always #(CFG_AVMM_CLK_PERIOD/2) i_cfg_avmm_clk = ~i_cfg_avmm_clk;
      always #(OSC_CLK_PERIOD/2)      i_osc_clk      = ~i_osc_clk;
      always #(PMA_CLK_PERIOD/2)      i_rx_pma_clk   = ~i_rx_pma_clk;
      always #(PMA_CLK_PERIOD)        i_rx_pma_div2_clk = ~i_rx_pma_div2_clk;
      always #(PMA_CLK_PERIOD/2)      i_tx_pma_clk   = ~i_tx_pma_clk;

     //=================================================================================
    //Below are DFx related signals, temporarily tie them off to 0s, need to be changed later
    logic i_scan_clk,
          i_test_clk_125m,
          i_test_clk_1g,
          i_test_clk_250m,
          i_test_clk_500m,
          i_test_clk_62m;

    logic [`AIBADAPTWRAPTCB_SCAN_CHAINS_RNG] i_test_c3adapt_scan_in;
    logic [`AIBADAPTWRAPTCB_STATIC_COMMON_RNG] i_test_c3adapt_tcb_static_common;
    logic [`AIBADAPTWRAPTCB_SCAN_CHAINS_RNG]   o_test_c3adapt_scan_out;
    logic [`AIBADAPTWRAPTCB_JTAG_OUT_RNG]      o_test_c3adapttcb_jtag;
    
    logic i_jtag_rstb_in,
          i_jtag_rstb_en_in,
          i_jtag_clkdr_in,
          i_jtag_clksel_in,
          i_jtag_intest_in,
          i_jtag_mode_in,
          i_jtag_weakpdn_in,
          i_jtag_weakpu_in,
          i_jtag_bs_scanen_in,
          i_jtag_bs_chain_in,
          i_jtag_last_bs_chain_in,
          i_por_aib_vcchssi,
          i_por_aib_vccl,
          i_red_idataselb_in_chain1,
          i_red_idataselb_in_chain2,
          i_red_shift_en_in_chain1,
          i_red_shift_en_in_chain2,
          i_txen_in_chain1,
          i_txen_in_chain2,
          i_directout_data_chain1_in,
          i_directout_data_chain2_in;

    initial begin
        i_scan_clk      = 1'b0;
        i_test_clk_125m = 1'b0;
        i_test_clk_1g   = 1'b0;
        i_test_clk_250m = 1'b0;
        i_test_clk_500m = 1'b0;
        i_test_clk_62m  = 1'b0;

        i_jtag_rstb_in = 1'b0;
        i_jtag_rstb_en_in = 1'b0;
        i_jtag_clkdr_in = 1'b0;
        i_jtag_clksel_in = 1'b0;
        i_jtag_intest_in = 1'b0;
        i_jtag_mode_in = 1'b0;
        i_jtag_weakpdn_in = 1'b0;
        i_jtag_weakpu_in = 1'b0;
        i_jtag_bs_scanen_in = 1'b0;
        i_jtag_bs_chain_in = 1'b0;
        i_jtag_last_bs_chain_in = 0;
        i_por_aib_vcchssi = 1'b0;
        i_por_aib_vccl = 1'b0;
        i_red_idataselb_in_chain1 = 1'b0;
        i_red_idataselb_in_chain2 = 1'b0;
        i_red_shift_en_in_chain1 = 1'b0;
        i_red_shift_en_in_chain2 = 1'b0;
        i_txen_in_chain1 = 1'b0;
        i_txen_in_chain2 = 1'b0;
        i_directout_data_chain1_in = 1'b0;
        i_directout_data_chain2_in = 1'b0;
        i_test_c3adapt_scan_in = 0;
        i_test_c3adapt_tcb_static_common = 0;
                
    end // initial begin

    //=================================================================================
    // AIB IOs
/*
    wire      aib0; 
    wire      aib1; 
    wire      aib10;
    wire      aib11;
    wire      aib12;
    wire      aib13;
    wire      aib14;
    wire      aib15;
    wire      aib16;
    wire      aib17;
    wire      aib18;
    wire      aib19;
    wire      aib2; 
    wire      aib20;
    wire      aib21;
    wire      aib22;
    wire      aib23;
    wire      aib24;
    wire      aib25;
    wire      aib26;
    wire      aib27;
    wire      aib28;
    wire      aib29;
    wire      aib3; 
    wire      aib30;
    wire      aib31;
    wire      aib32;
    wire      aib33;
    wire      aib34;
    wire      aib35;
    wire      aib36;
    wire      aib37;
    wire      aib38;
    wire      aib39;
    wire      aib4; 
    wire      aib40;
    wire      aib41;
    wire      aib42;
    wire      aib43;
    wire      aib44;
    wire      aib45;
    wire      aib46;
    wire      aib47;
    wire      aib48;
    wire      aib49;
    wire      aib5; 
    wire      aib50;
    wire      aib51;
    wire      aib52;
    wire      aib53;
    wire      aib54;
    wire      aib55;
    wire      aib56;
    wire      aib57;
    wire      aib58;
    wire      aib59;
    wire      aib6; 
    wire      aib60;
    wire      aib61;
    wire      aib62;
    wire      aib63;
    wire      aib64;
    wire      aib65;
    wire      aib66;
    wire      aib67;
    wire      aib68;
    wire      aib69;
    wire      aib7; 
    wire      aib70;
    wire      aib71;
    wire      aib72;
    wire      aib73;
    wire      aib74;
    wire      aib75;
    wire      aib76;
    wire      aib77;
    wire      aib78;
    wire      aib79;
    wire      aib8; 
    wire      aib80;
    wire      aib81;
    wire      aib82;
    wire      aib83;
    wire      aib84;
    wire      aib85;
    wire      aib86;
    wire      aib87;
    wire      aib88;
    wire      aib89;
    wire      aib9; 
    wire      aib90;
    wire      aib91;
    wire      aib92;
    wire      aib93;
    wire      aib94;
    wire      aib95;

    wire      aib20_o;
    wire      aib21_o;
    wire      aib22_o;
    wire      aib23_o;
    wire      aib24_o;
    wire      aib25_o;
    wire      aib26_o;
    wire      aib27_o;
    wire      aib28_o;
    wire      aib29_o;
    wire      aib30_o;
    wire      aib31_o;
    wire      aib32_o;
    wire      aib33_o;
    wire      aib34_o;
    wire      aib35_o;
    wire      aib36_o;
    wire      aib37_o;
    wire      aib38_o;
    wire      aib39_o;

    wire      aib40_o;
    wire      aib41_o;
    wire      aib82_o;
    wire      aib83_o;
 */   
    /*AUTOWIRE*/
    // Beginning of automatic wires (for undeclared instantiated-module outputs)
    wire [16:0]         o_adpt_cfg_addr;        // From dut of c3aibadapt_wrap.v
    wire [3:0]          o_adpt_cfg_byte_en;     // From dut of c3aibadapt_wrap.v
    wire                o_adpt_cfg_clk;         // From dut of c3aibadapt_wrap.v
    wire                o_adpt_cfg_read;        // From dut of c3aibadapt_wrap.v
    wire                o_adpt_cfg_rst_n;       // From dut of c3aibadapt_wrap.v
    wire [31:0]         o_adpt_cfg_wdata;       // From dut of c3aibadapt_wrap.v
    wire                o_adpt_cfg_write;       // From dut of c3aibadapt_wrap.v
    wire                o_adpt_hard_rst_n;      // From dut of c3aibadapt_wrap.v
    wire [12:0]         o_aibdftdll2adjch;      // From dut of c3aibadapt_wrap.v
    wire [31:0]         o_cfg_avmm_rdata;       // From dut of c3aibadapt_wrap.v
    wire                o_cfg_avmm_rdatavld;    // From dut of c3aibadapt_wrap.v
    wire                o_cfg_avmm_waitreq;     // From dut of c3aibadapt_wrap.v
    wire [60:0]         o_chnl_ssr;             // From dut of c3aibadapt_wrap.v
    wire                o_directout_data_chain1_out;// From dut of c3aibadapt_wrap.v
    wire                o_directout_data_chain2_out;// From dut of c3aibadapt_wrap.v
    wire [2:0]          o_ehip_init_status;     // From dut of c3aibadapt_wrap.v
    wire                o_jtag_bs_chain_out;    // From dut of c3aibadapt_wrap.v
    wire                o_jtag_bs_scanen_out;   // From dut of c3aibadapt_wrap.v
    wire                o_jtag_clkdr_out;       // From dut of c3aibadapt_wrap.v
    wire                o_jtag_clksel_out;      // From dut of c3aibadapt_wrap.v
    wire                o_jtag_intest_out;      // From dut of c3aibadapt_wrap.v
    wire                o_jtag_last_bs_chain_out;// From dut of c3aibadapt_wrap.v
    wire                o_jtag_mode_out;        // From dut of c3aibadapt_wrap.v
    wire                o_jtag_rstb_en_out;     // From dut of c3aibadapt_wrap.v
    wire                o_jtag_rstb_out;        // From dut of c3aibadapt_wrap.v
    wire                o_jtag_weakpdn_out;     // From dut of c3aibadapt_wrap.v
    wire                o_jtag_weakpu_out;      // From dut of c3aibadapt_wrap.v
    wire                o_osc_clk;              // From dut of c3aibadapt_wrap.v
    wire                o_por_aib_vcchssi;      // From dut of c3aibadapt_wrap.v
    wire                o_por_aib_vccl;         // From dut of c3aibadapt_wrap.v
    wire                o_red_idataselb_out_chain1;// From dut of c3aibadapt_wrap.v
    wire                o_red_idataselb_out_chain2;// From dut of c3aibadapt_wrap.v
    wire                o_red_shift_en_out_chain1;// From dut of c3aibadapt_wrap.v
    wire                o_red_shift_en_out_chain2;// From dut of c3aibadapt_wrap.v
    wire                o_rx_xcvrif_rst_n;      // From dut of c3aibadapt_wrap.v
//  wire [39:0]         o_tx_pma_data;          // From dut of c3aibadapt_wrap.v
    wire                o_tx_transfer_clk;      // From dut of c3aibadapt_wrap.v
    logic [23:0]        o_tx_transfer_div2_clk; // From dut of c3aibadapt_wrap.v
    wire                o_tx_xcvrif_rst_n;      // From dut of c3aibadapt_wrap.v
    wire                o_txen_out_chain1;      // From dut of c3aibadapt_wrap.v
    wire                o_txen_out_chain2;      // From dut of c3aibadapt_wrap.v
    wire                HI;
    wire                LO;
    wire  [81*24-1:0]   ms_sideband;
    wire  [73*24-1:0]   sl_sideband;              
    // End of automatics
   // EMIB Side
// wire [95:0] AIB_CHAN0;
   wire [95:0] AIB_CHAN1;
   wire [95:0] AIB_CHAN2;
   wire [95:0] AIB_CHAN3;
   wire [95:0] AIB_CHAN4;
   wire [95:0] AIB_CHAN5;
   wire [95:0] AIB_CHAN6;
   wire [95:0] AIB_CHAN7;
   wire [95:0] AIB_CHAN8;
   wire [95:0] AIB_CHAN9;
   wire [95:0] AIB_CHAN10;
   wire [95:0] AIB_CHAN11;
   wire [95:0] AIB_CHAN12;
   wire [95:0] AIB_CHAN13;
   wire [95:0] AIB_CHAN14;
   wire [95:0] AIB_CHAN15;
   wire [95:0] AIB_CHAN16;
   wire [95:0] AIB_CHAN17;
   wire [95:0] AIB_CHAN18;
   wire [95:0] AIB_CHAN19;
   wire [95:0] AIB_CHAN20;
   wire [95:0] AIB_CHAN21;
   wire [95:0] AIB_CHAN22;
   wire [95:0] AIB_CHAN23;
   wire [95:0] AIB_AUX;
/*
    wire        aib95_ch0_x0y0, aib94_ch0_x0y0, aib93_ch0_x0y0,aib92_ch0_x0y0,
                aib91_ch0_x0y0, aib90_ch0_x0y0, aib89_ch0_x0y0,aib88_ch0_x0y0,
                aib87_ch0_x0y0, aib86_ch0_x0y0, aib85_ch0_x0y0,aib84_ch0_x0y0,
                aib83_ch0_x0y0, aib82_ch0_x0y0, aib81_ch0_x0y0,aib80_ch0_x0y0,
                aib79_ch0_x0y0, aib78_ch0_x0y0, aib77_ch0_x0y0,aib76_ch0_x0y0,
                aib75_ch0_x0y0, aib74_ch0_x0y0, aib73_ch0_x0y0,aib72_ch0_x0y0,
                aib71_ch0_x0y0, aib70_ch0_x0y0, aib69_ch0_x0y0,aib68_ch0_x0y0,
                aib67_ch0_x0y0, aib66_ch0_x0y0, aib65_ch0_x0y0,aib64_ch0_x0y0,
                aib63_ch0_x0y0, aib62_ch0_x0y0, aib61_ch0_x0y0,aib60_ch0_x0y0,
                aib59_ch0_x0y0, aib58_ch0_x0y0, aib57_ch0_x0y0,aib56_ch0_x0y0,
                aib55_ch0_x0y0, aib54_ch0_x0y0, aib53_ch0_x0y0,aib52_ch0_x0y0,
                aib51_ch0_x0y0, aib50_ch0_x0y0, aib49_ch0_x0y0,aib48_ch0_x0y0,
                aib47_ch0_x0y0, aib46_ch0_x0y0, aib45_ch0_x0y0,aib44_ch0_x0y0,
                aib43_ch0_x0y0, aib42_ch0_x0y0, aib41_ch0_x0y0,aib40_ch0_x0y0,
                aib39_ch0_x0y0, aib38_ch0_x0y0, aib37_ch0_x0y0,aib36_ch0_x0y0,
                aib35_ch0_x0y0, aib34_ch0_x0y0, aib33_ch0_x0y0,aib32_ch0_x0y0,
                aib31_ch0_x0y0, aib30_ch0_x0y0, aib29_ch0_x0y0,aib28_ch0_x0y0,
                aib27_ch0_x0y0, aib26_ch0_x0y0, aib25_ch0_x0y0,aib24_ch0_x0y0,
                aib23_ch0_x0y0, aib22_ch0_x0y0, aib21_ch0_x0y0,aib20_ch0_x0y0,
                aib19_ch0_x0y0, aib18_ch0_x0y0, aib17_ch0_x0y0,aib16_ch0_x0y0,
                aib15_ch0_x0y0, aib14_ch0_x0y0, aib13_ch0_x0y0,aib12_ch0_x0y0,
                aib11_ch0_x0y0, aib10_ch0_x0y0, aib9_ch0_x0y0,aib8_ch0_x0y0,
                aib7_ch0_x0y0, aib6_ch0_x0y0, aib5_ch0_x0y0,aib4_ch0_x0y0,
                aib3_ch0_x0y0, aib2_ch0_x0y0, aib1_ch0_x0y0,aib0_ch0_x0y0;
    assign aib82_ch0_x0y0 = aib84_ch0_x0y0;
    assign aib83_ch0_x0y0 = aib85_ch0_x0y0;
*/
    wire        aib95_ch1_x0y0, aib94_ch1_x0y0, aib93_ch1_x0y0,aib92_ch1_x0y0,
                aib91_ch1_x0y0, aib90_ch1_x0y0, aib89_ch1_x0y0,aib88_ch1_x0y0,
                aib87_ch1_x0y0, aib86_ch1_x0y0, aib85_ch1_x0y0,aib84_ch1_x0y0,
                aib83_ch1_x0y0, aib82_ch1_x0y0, aib81_ch1_x0y0,aib80_ch1_x0y0,
                aib79_ch1_x0y0, aib78_ch1_x0y0, aib77_ch1_x0y0,aib76_ch1_x0y0,
                aib75_ch1_x0y0, aib74_ch1_x0y0, aib73_ch1_x0y0,aib72_ch1_x0y0,
                aib71_ch1_x0y0, aib70_ch1_x0y0, aib69_ch1_x0y0,aib68_ch1_x0y0,
                aib67_ch1_x0y0, aib66_ch1_x0y0, aib65_ch1_x0y0,aib64_ch1_x0y0,
                aib63_ch1_x0y0, aib62_ch1_x0y0, aib61_ch1_x0y0,aib60_ch1_x0y0,
                aib59_ch1_x0y0, aib58_ch1_x0y0, aib57_ch1_x0y0,aib56_ch1_x0y0,
                aib55_ch1_x0y0, aib54_ch1_x0y0, aib53_ch1_x0y0,aib52_ch1_x0y0,
                aib51_ch1_x0y0, aib50_ch1_x0y0, aib49_ch1_x0y0,aib48_ch1_x0y0,
                aib47_ch1_x0y0, aib46_ch1_x0y0, aib45_ch1_x0y0,aib44_ch1_x0y0,
                aib43_ch1_x0y0, aib42_ch1_x0y0, aib41_ch1_x0y0,aib40_ch1_x0y0,
                aib39_ch1_x0y0, aib38_ch1_x0y0, aib37_ch1_x0y0,aib36_ch1_x0y0,
                aib35_ch1_x0y0, aib34_ch1_x0y0, aib33_ch1_x0y0,aib32_ch1_x0y0,
                aib31_ch1_x0y0, aib30_ch1_x0y0, aib29_ch1_x0y0,aib28_ch1_x0y0,
                aib27_ch1_x0y0, aib26_ch1_x0y0, aib25_ch1_x0y0,aib24_ch1_x0y0,
                aib23_ch1_x0y0, aib22_ch1_x0y0, aib21_ch1_x0y0,aib20_ch1_x0y0,
                aib19_ch1_x0y0, aib18_ch1_x0y0, aib17_ch1_x0y0,aib16_ch1_x0y0,
                aib15_ch1_x0y0, aib14_ch1_x0y0, aib13_ch1_x0y0,aib12_ch1_x0y0,
                aib11_ch1_x0y0, aib10_ch1_x0y0, aib9_ch1_x0y0,aib8_ch1_x0y0,
                aib7_ch1_x0y0, aib6_ch1_x0y0, aib5_ch1_x0y0,aib4_ch1_x0y0,
                aib3_ch1_x0y0, aib2_ch1_x0y0, aib1_ch1_x0y0,aib0_ch1_x0y0;
    wire        aib95_ch2_x0y0, aib94_ch2_x0y0, aib93_ch2_x0y0,aib92_ch2_x0y0,
                aib91_ch2_x0y0, aib90_ch2_x0y0, aib89_ch2_x0y0,aib88_ch2_x0y0,
                aib87_ch2_x0y0, aib86_ch2_x0y0, aib85_ch2_x0y0,aib84_ch2_x0y0,
                aib83_ch2_x0y0, aib82_ch2_x0y0, aib81_ch2_x0y0,aib80_ch2_x0y0,
                aib79_ch2_x0y0, aib78_ch2_x0y0, aib77_ch2_x0y0,aib76_ch2_x0y0,
                aib75_ch2_x0y0, aib74_ch2_x0y0, aib73_ch2_x0y0,aib72_ch2_x0y0,
                aib71_ch2_x0y0, aib70_ch2_x0y0, aib69_ch2_x0y0,aib68_ch2_x0y0,
                aib67_ch2_x0y0, aib66_ch2_x0y0, aib65_ch2_x0y0,aib64_ch2_x0y0,
                aib63_ch2_x0y0, aib62_ch2_x0y0, aib61_ch2_x0y0,aib60_ch2_x0y0,
                aib59_ch2_x0y0, aib58_ch2_x0y0, aib57_ch2_x0y0,aib56_ch2_x0y0,
                aib55_ch2_x0y0, aib54_ch2_x0y0, aib53_ch2_x0y0,aib52_ch2_x0y0,
                aib51_ch2_x0y0, aib50_ch2_x0y0, aib49_ch2_x0y0,aib48_ch2_x0y0,
                aib47_ch2_x0y0, aib46_ch2_x0y0, aib45_ch2_x0y0,aib44_ch2_x0y0,
                aib43_ch2_x0y0, aib42_ch2_x0y0, aib41_ch2_x0y0,aib40_ch2_x0y0,
                aib39_ch2_x0y0, aib38_ch2_x0y0, aib37_ch2_x0y0,aib36_ch2_x0y0,
                aib35_ch2_x0y0, aib34_ch2_x0y0, aib33_ch2_x0y0,aib32_ch2_x0y0,
                aib31_ch2_x0y0, aib30_ch2_x0y0, aib29_ch2_x0y0,aib28_ch2_x0y0,
                aib27_ch2_x0y0, aib26_ch2_x0y0, aib25_ch2_x0y0,aib24_ch2_x0y0,
                aib23_ch2_x0y0, aib22_ch2_x0y0, aib21_ch2_x0y0,aib20_ch2_x0y0,
                aib19_ch2_x0y0, aib18_ch2_x0y0, aib17_ch2_x0y0,aib16_ch2_x0y0,
                aib15_ch2_x0y0, aib14_ch2_x0y0, aib13_ch2_x0y0,aib12_ch2_x0y0,
                aib11_ch2_x0y0, aib10_ch2_x0y0, aib9_ch2_x0y0,aib8_ch2_x0y0,
                aib7_ch2_x0y0, aib6_ch2_x0y0, aib5_ch2_x0y0,aib4_ch2_x0y0,
                aib3_ch2_x0y0, aib2_ch2_x0y0, aib1_ch2_x0y0,aib0_ch2_x0y0; 
    wire        aib95_ch3_x0y0, aib94_ch3_x0y0, aib93_ch3_x0y0,aib92_ch3_x0y0,
                aib91_ch3_x0y0, aib90_ch3_x0y0, aib89_ch3_x0y0,aib88_ch3_x0y0,
                aib87_ch3_x0y0, aib86_ch3_x0y0, aib85_ch3_x0y0,aib84_ch3_x0y0,
                aib83_ch3_x0y0, aib82_ch3_x0y0, aib81_ch3_x0y0,aib80_ch3_x0y0,
                aib79_ch3_x0y0, aib78_ch3_x0y0, aib77_ch3_x0y0,aib76_ch3_x0y0,
                aib75_ch3_x0y0, aib74_ch3_x0y0, aib73_ch3_x0y0,aib72_ch3_x0y0,
                aib71_ch3_x0y0, aib70_ch3_x0y0, aib69_ch3_x0y0,aib68_ch3_x0y0,
                aib67_ch3_x0y0, aib66_ch3_x0y0, aib65_ch3_x0y0,aib64_ch3_x0y0,
                aib63_ch3_x0y0, aib62_ch3_x0y0, aib61_ch3_x0y0,aib60_ch3_x0y0,
                aib59_ch3_x0y0, aib58_ch3_x0y0, aib57_ch3_x0y0,aib56_ch3_x0y0,
                aib55_ch3_x0y0, aib54_ch3_x0y0, aib53_ch3_x0y0,aib52_ch3_x0y0,
                aib51_ch3_x0y0, aib50_ch3_x0y0, aib49_ch3_x0y0,aib48_ch3_x0y0,
                aib47_ch3_x0y0, aib46_ch3_x0y0, aib45_ch3_x0y0,aib44_ch3_x0y0,
                aib43_ch3_x0y0, aib42_ch3_x0y0, aib41_ch3_x0y0,aib40_ch3_x0y0,
                aib39_ch3_x0y0, aib38_ch3_x0y0, aib37_ch3_x0y0,aib36_ch3_x0y0,
                aib35_ch3_x0y0, aib34_ch3_x0y0, aib33_ch3_x0y0,aib32_ch3_x0y0,
                aib31_ch3_x0y0, aib30_ch3_x0y0, aib29_ch3_x0y0,aib28_ch3_x0y0,
                aib27_ch3_x0y0, aib26_ch3_x0y0, aib25_ch3_x0y0,aib24_ch3_x0y0,
                aib23_ch3_x0y0, aib22_ch3_x0y0, aib21_ch3_x0y0,aib20_ch3_x0y0,
                aib19_ch3_x0y0, aib18_ch3_x0y0, aib17_ch3_x0y0,aib16_ch3_x0y0,
                aib15_ch3_x0y0, aib14_ch3_x0y0, aib13_ch3_x0y0,aib12_ch3_x0y0,
                aib11_ch3_x0y0, aib10_ch3_x0y0, aib9_ch3_x0y0,aib8_ch3_x0y0,
                aib7_ch3_x0y0, aib6_ch3_x0y0, aib5_ch3_x0y0,aib4_ch3_x0y0,
                aib3_ch3_x0y0, aib2_ch3_x0y0, aib1_ch3_x0y0,aib0_ch3_x0y0;
    wire        aib95_ch4_x0y0, aib94_ch4_x0y0, aib93_ch4_x0y0,aib92_ch4_x0y0,
                aib91_ch4_x0y0, aib90_ch4_x0y0, aib89_ch4_x0y0,aib88_ch4_x0y0,
                aib87_ch4_x0y0, aib86_ch4_x0y0, aib85_ch4_x0y0,aib84_ch4_x0y0,
                aib83_ch4_x0y0, aib82_ch4_x0y0, aib81_ch4_x0y0,aib80_ch4_x0y0,
                aib79_ch4_x0y0, aib78_ch4_x0y0, aib77_ch4_x0y0,aib76_ch4_x0y0,
                aib75_ch4_x0y0, aib74_ch4_x0y0, aib73_ch4_x0y0,aib72_ch4_x0y0,
                aib71_ch4_x0y0, aib70_ch4_x0y0, aib69_ch4_x0y0,aib68_ch4_x0y0,
                aib67_ch4_x0y0, aib66_ch4_x0y0, aib65_ch4_x0y0,aib64_ch4_x0y0,
                aib63_ch4_x0y0, aib62_ch4_x0y0, aib61_ch4_x0y0,aib60_ch4_x0y0,
                aib59_ch4_x0y0, aib58_ch4_x0y0, aib57_ch4_x0y0,aib56_ch4_x0y0,
                aib55_ch4_x0y0, aib54_ch4_x0y0, aib53_ch4_x0y0,aib52_ch4_x0y0,
                aib51_ch4_x0y0, aib50_ch4_x0y0, aib49_ch4_x0y0,aib48_ch4_x0y0,
                aib47_ch4_x0y0, aib46_ch4_x0y0, aib45_ch4_x0y0,aib44_ch4_x0y0,
                aib43_ch4_x0y0, aib42_ch4_x0y0, aib41_ch4_x0y0,aib40_ch4_x0y0,
                aib39_ch4_x0y0, aib38_ch4_x0y0, aib37_ch4_x0y0,aib36_ch4_x0y0,
                aib35_ch4_x0y0, aib34_ch4_x0y0, aib33_ch4_x0y0,aib32_ch4_x0y0,
                aib31_ch4_x0y0, aib30_ch4_x0y0, aib29_ch4_x0y0,aib28_ch4_x0y0,
                aib27_ch4_x0y0, aib26_ch4_x0y0, aib25_ch4_x0y0,aib24_ch4_x0y0,
                aib23_ch4_x0y0, aib22_ch4_x0y0, aib21_ch4_x0y0,aib20_ch4_x0y0,
                aib19_ch4_x0y0, aib18_ch4_x0y0, aib17_ch4_x0y0,aib16_ch4_x0y0,
                aib15_ch4_x0y0, aib14_ch4_x0y0, aib13_ch4_x0y0,aib12_ch4_x0y0,
                aib11_ch4_x0y0, aib10_ch4_x0y0, aib9_ch4_x0y0,aib8_ch4_x0y0,
                aib7_ch4_x0y0, aib6_ch4_x0y0, aib5_ch4_x0y0,aib4_ch4_x0y0,
                aib3_ch4_x0y0, aib2_ch4_x0y0, aib1_ch4_x0y0,aib0_ch4_x0y0; 
    wire        aib95_ch5_x0y0, aib94_ch5_x0y0, aib93_ch5_x0y0,aib92_ch5_x0y0,
                aib91_ch5_x0y0, aib90_ch5_x0y0, aib89_ch5_x0y0,aib88_ch5_x0y0,
                aib87_ch5_x0y0, aib86_ch5_x0y0, aib85_ch5_x0y0,aib84_ch5_x0y0,
                aib83_ch5_x0y0, aib82_ch5_x0y0, aib81_ch5_x0y0,aib80_ch5_x0y0,
                aib79_ch5_x0y0, aib78_ch5_x0y0, aib77_ch5_x0y0,aib76_ch5_x0y0,
                aib75_ch5_x0y0, aib74_ch5_x0y0, aib73_ch5_x0y0,aib72_ch5_x0y0,
                aib71_ch5_x0y0, aib70_ch5_x0y0, aib69_ch5_x0y0,aib68_ch5_x0y0,
                aib67_ch5_x0y0, aib66_ch5_x0y0, aib65_ch5_x0y0,aib64_ch5_x0y0,
                aib63_ch5_x0y0, aib62_ch5_x0y0, aib61_ch5_x0y0,aib60_ch5_x0y0,
                aib59_ch5_x0y0, aib58_ch5_x0y0, aib57_ch5_x0y0,aib56_ch5_x0y0,
                aib55_ch5_x0y0, aib54_ch5_x0y0, aib53_ch5_x0y0,aib52_ch5_x0y0,
                aib51_ch5_x0y0, aib50_ch5_x0y0, aib49_ch5_x0y0,aib48_ch5_x0y0,
                aib47_ch5_x0y0, aib46_ch5_x0y0, aib45_ch5_x0y0,aib44_ch5_x0y0,
                aib43_ch5_x0y0, aib42_ch5_x0y0, aib41_ch5_x0y0,aib40_ch5_x0y0,
                aib39_ch5_x0y0, aib38_ch5_x0y0, aib37_ch5_x0y0,aib36_ch5_x0y0,
                aib35_ch5_x0y0, aib34_ch5_x0y0, aib33_ch5_x0y0,aib32_ch5_x0y0,
                aib31_ch5_x0y0, aib30_ch5_x0y0, aib29_ch5_x0y0,aib28_ch5_x0y0,
                aib27_ch5_x0y0, aib26_ch5_x0y0, aib25_ch5_x0y0,aib24_ch5_x0y0,
                aib23_ch5_x0y0, aib22_ch5_x0y0, aib21_ch5_x0y0,aib20_ch5_x0y0,
                aib19_ch5_x0y0, aib18_ch5_x0y0, aib17_ch5_x0y0,aib16_ch5_x0y0,
                aib15_ch5_x0y0, aib14_ch5_x0y0, aib13_ch5_x0y0,aib12_ch5_x0y0,
                aib11_ch5_x0y0, aib10_ch5_x0y0, aib9_ch5_x0y0,aib8_ch5_x0y0,
                aib7_ch5_x0y0, aib6_ch5_x0y0, aib5_ch5_x0y0,aib4_ch5_x0y0,
                aib3_ch5_x0y0, aib2_ch5_x0y0, aib1_ch5_x0y0,aib0_ch5_x0y0;
    wire        aib95_ch0_x0y1, aib94_ch0_x0y1, aib93_ch0_x0y1,aib92_ch0_x0y1,
                aib91_ch0_x0y1, aib90_ch0_x0y1, aib89_ch0_x0y1,aib88_ch0_x0y1,
                aib87_ch0_x0y1, aib86_ch0_x0y1, aib85_ch0_x0y1,aib84_ch0_x0y1,
                aib83_ch0_x0y1, aib82_ch0_x0y1, aib81_ch0_x0y1,aib80_ch0_x0y1,
                aib79_ch0_x0y1, aib78_ch0_x0y1, aib77_ch0_x0y1,aib76_ch0_x0y1,
                aib75_ch0_x0y1, aib74_ch0_x0y1, aib73_ch0_x0y1,aib72_ch0_x0y1,
                aib71_ch0_x0y1, aib70_ch0_x0y1, aib69_ch0_x0y1,aib68_ch0_x0y1,
                aib67_ch0_x0y1, aib66_ch0_x0y1, aib65_ch0_x0y1,aib64_ch0_x0y1,
                aib63_ch0_x0y1, aib62_ch0_x0y1, aib61_ch0_x0y1,aib60_ch0_x0y1,
                aib59_ch0_x0y1, aib58_ch0_x0y1, aib57_ch0_x0y1,aib56_ch0_x0y1,
                aib55_ch0_x0y1, aib54_ch0_x0y1, aib53_ch0_x0y1,aib52_ch0_x0y1,
                aib51_ch0_x0y1, aib50_ch0_x0y1, aib49_ch0_x0y1,aib48_ch0_x0y1,
                aib47_ch0_x0y1, aib46_ch0_x0y1, aib45_ch0_x0y1,aib44_ch0_x0y1,
                aib43_ch0_x0y1, aib42_ch0_x0y1, aib41_ch0_x0y1,aib40_ch0_x0y1,
                aib39_ch0_x0y1, aib38_ch0_x0y1, aib37_ch0_x0y1,aib36_ch0_x0y1,
                aib35_ch0_x0y1, aib34_ch0_x0y1, aib33_ch0_x0y1,aib32_ch0_x0y1,
                aib31_ch0_x0y1, aib30_ch0_x0y1, aib29_ch0_x0y1,aib28_ch0_x0y1,
                aib27_ch0_x0y1, aib26_ch0_x0y1, aib25_ch0_x0y1,aib24_ch0_x0y1,
                aib23_ch0_x0y1, aib22_ch0_x0y1, aib21_ch0_x0y1,aib20_ch0_x0y1,
                aib19_ch0_x0y1, aib18_ch0_x0y1, aib17_ch0_x0y1,aib16_ch0_x0y1,
                aib15_ch0_x0y1, aib14_ch0_x0y1, aib13_ch0_x0y1,aib12_ch0_x0y1,
                aib11_ch0_x0y1, aib10_ch0_x0y1, aib9_ch0_x0y1,aib8_ch0_x0y1,
                aib7_ch0_x0y1, aib6_ch0_x0y1, aib5_ch0_x0y1,aib4_ch0_x0y1,
                aib3_ch0_x0y1, aib2_ch0_x0y1, aib1_ch0_x0y1,aib0_ch0_x0y1;
    wire        aib95_ch1_x0y1, aib94_ch1_x0y1, aib93_ch1_x0y1,aib92_ch1_x0y1,
                aib91_ch1_x0y1, aib90_ch1_x0y1, aib89_ch1_x0y1,aib88_ch1_x0y1,
                aib87_ch1_x0y1, aib86_ch1_x0y1, aib85_ch1_x0y1,aib84_ch1_x0y1,
                aib83_ch1_x0y1, aib82_ch1_x0y1, aib81_ch1_x0y1,aib80_ch1_x0y1,
                aib79_ch1_x0y1, aib78_ch1_x0y1, aib77_ch1_x0y1,aib76_ch1_x0y1,
                aib75_ch1_x0y1, aib74_ch1_x0y1, aib73_ch1_x0y1,aib72_ch1_x0y1,
                aib71_ch1_x0y1, aib70_ch1_x0y1, aib69_ch1_x0y1,aib68_ch1_x0y1,
                aib67_ch1_x0y1, aib66_ch1_x0y1, aib65_ch1_x0y1,aib64_ch1_x0y1,
                aib63_ch1_x0y1, aib62_ch1_x0y1, aib61_ch1_x0y1,aib60_ch1_x0y1,
                aib59_ch1_x0y1, aib58_ch1_x0y1, aib57_ch1_x0y1,aib56_ch1_x0y1,
                aib55_ch1_x0y1, aib54_ch1_x0y1, aib53_ch1_x0y1,aib52_ch1_x0y1,
                aib51_ch1_x0y1, aib50_ch1_x0y1, aib49_ch1_x0y1,aib48_ch1_x0y1,
                aib47_ch1_x0y1, aib46_ch1_x0y1, aib45_ch1_x0y1,aib44_ch1_x0y1,
                aib43_ch1_x0y1, aib42_ch1_x0y1, aib41_ch1_x0y1,aib40_ch1_x0y1,
                aib39_ch1_x0y1, aib38_ch1_x0y1, aib37_ch1_x0y1,aib36_ch1_x0y1,
                aib35_ch1_x0y1, aib34_ch1_x0y1, aib33_ch1_x0y1,aib32_ch1_x0y1,
                aib31_ch1_x0y1, aib30_ch1_x0y1, aib29_ch1_x0y1,aib28_ch1_x0y1,
                aib27_ch1_x0y1, aib26_ch1_x0y1, aib25_ch1_x0y1,aib24_ch1_x0y1,
                aib23_ch1_x0y1, aib22_ch1_x0y1, aib21_ch1_x0y1,aib20_ch1_x0y1,
                aib19_ch1_x0y1, aib18_ch1_x0y1, aib17_ch1_x0y1,aib16_ch1_x0y1,
                aib15_ch1_x0y1, aib14_ch1_x0y1, aib13_ch1_x0y1,aib12_ch1_x0y1,
                aib11_ch1_x0y1, aib10_ch1_x0y1, aib9_ch1_x0y1,aib8_ch1_x0y1,
                aib7_ch1_x0y1, aib6_ch1_x0y1, aib5_ch1_x0y1,aib4_ch1_x0y1,
                aib3_ch1_x0y1, aib2_ch1_x0y1, aib1_ch1_x0y1,aib0_ch1_x0y1;
    wire        aib95_ch2_x0y1, aib94_ch2_x0y1, aib93_ch2_x0y1,aib92_ch2_x0y1,
                aib91_ch2_x0y1, aib90_ch2_x0y1, aib89_ch2_x0y1,aib88_ch2_x0y1,
                aib87_ch2_x0y1, aib86_ch2_x0y1, aib85_ch2_x0y1,aib84_ch2_x0y1,
                aib83_ch2_x0y1, aib82_ch2_x0y1, aib81_ch2_x0y1,aib80_ch2_x0y1,
                aib79_ch2_x0y1, aib78_ch2_x0y1, aib77_ch2_x0y1,aib76_ch2_x0y1,
                aib75_ch2_x0y1, aib74_ch2_x0y1, aib73_ch2_x0y1,aib72_ch2_x0y1,
                aib71_ch2_x0y1, aib70_ch2_x0y1, aib69_ch2_x0y1,aib68_ch2_x0y1,
                aib67_ch2_x0y1, aib66_ch2_x0y1, aib65_ch2_x0y1,aib64_ch2_x0y1,
                aib63_ch2_x0y1, aib62_ch2_x0y1, aib61_ch2_x0y1,aib60_ch2_x0y1,
                aib59_ch2_x0y1, aib58_ch2_x0y1, aib57_ch2_x0y1,aib56_ch2_x0y1,
                aib55_ch2_x0y1, aib54_ch2_x0y1, aib53_ch2_x0y1,aib52_ch2_x0y1,
                aib51_ch2_x0y1, aib50_ch2_x0y1, aib49_ch2_x0y1,aib48_ch2_x0y1,
                aib47_ch2_x0y1, aib46_ch2_x0y1, aib45_ch2_x0y1,aib44_ch2_x0y1,
                aib43_ch2_x0y1, aib42_ch2_x0y1, aib41_ch2_x0y1,aib40_ch2_x0y1,
                aib39_ch2_x0y1, aib38_ch2_x0y1, aib37_ch2_x0y1,aib36_ch2_x0y1,
                aib35_ch2_x0y1, aib34_ch2_x0y1, aib33_ch2_x0y1,aib32_ch2_x0y1,
                aib31_ch2_x0y1, aib30_ch2_x0y1, aib29_ch2_x0y1,aib28_ch2_x0y1,
                aib27_ch2_x0y1, aib26_ch2_x0y1, aib25_ch2_x0y1,aib24_ch2_x0y1,
                aib23_ch2_x0y1, aib22_ch2_x0y1, aib21_ch2_x0y1,aib20_ch2_x0y1,
                aib19_ch2_x0y1, aib18_ch2_x0y1, aib17_ch2_x0y1,aib16_ch2_x0y1,
                aib15_ch2_x0y1, aib14_ch2_x0y1, aib13_ch2_x0y1,aib12_ch2_x0y1,
                aib11_ch2_x0y1, aib10_ch2_x0y1, aib9_ch2_x0y1,aib8_ch2_x0y1,
                aib7_ch2_x0y1, aib6_ch2_x0y1, aib5_ch2_x0y1,aib4_ch2_x0y1,
                aib3_ch2_x0y1, aib2_ch2_x0y1, aib1_ch2_x0y1,aib0_ch2_x0y1; 
    wire        aib95_ch3_x0y1, aib94_ch3_x0y1, aib93_ch3_x0y1,aib92_ch3_x0y1,
                aib91_ch3_x0y1, aib90_ch3_x0y1, aib89_ch3_x0y1,aib88_ch3_x0y1,
                aib87_ch3_x0y1, aib86_ch3_x0y1, aib85_ch3_x0y1,aib84_ch3_x0y1,
                aib83_ch3_x0y1, aib82_ch3_x0y1, aib81_ch3_x0y1,aib80_ch3_x0y1,
                aib79_ch3_x0y1, aib78_ch3_x0y1, aib77_ch3_x0y1,aib76_ch3_x0y1,
                aib75_ch3_x0y1, aib74_ch3_x0y1, aib73_ch3_x0y1,aib72_ch3_x0y1,
                aib71_ch3_x0y1, aib70_ch3_x0y1, aib69_ch3_x0y1,aib68_ch3_x0y1,
                aib67_ch3_x0y1, aib66_ch3_x0y1, aib65_ch3_x0y1,aib64_ch3_x0y1,
                aib63_ch3_x0y1, aib62_ch3_x0y1, aib61_ch3_x0y1,aib60_ch3_x0y1,
                aib59_ch3_x0y1, aib58_ch3_x0y1, aib57_ch3_x0y1,aib56_ch3_x0y1,
                aib55_ch3_x0y1, aib54_ch3_x0y1, aib53_ch3_x0y1,aib52_ch3_x0y1,
                aib51_ch3_x0y1, aib50_ch3_x0y1, aib49_ch3_x0y1,aib48_ch3_x0y1,
                aib47_ch3_x0y1, aib46_ch3_x0y1, aib45_ch3_x0y1,aib44_ch3_x0y1,
                aib43_ch3_x0y1, aib42_ch3_x0y1, aib41_ch3_x0y1,aib40_ch3_x0y1,
                aib39_ch3_x0y1, aib38_ch3_x0y1, aib37_ch3_x0y1,aib36_ch3_x0y1,
                aib35_ch3_x0y1, aib34_ch3_x0y1, aib33_ch3_x0y1,aib32_ch3_x0y1,
                aib31_ch3_x0y1, aib30_ch3_x0y1, aib29_ch3_x0y1,aib28_ch3_x0y1,
                aib27_ch3_x0y1, aib26_ch3_x0y1, aib25_ch3_x0y1,aib24_ch3_x0y1,
                aib23_ch3_x0y1, aib22_ch3_x0y1, aib21_ch3_x0y1,aib20_ch3_x0y1,
                aib19_ch3_x0y1, aib18_ch3_x0y1, aib17_ch3_x0y1,aib16_ch3_x0y1,
                aib15_ch3_x0y1, aib14_ch3_x0y1, aib13_ch3_x0y1,aib12_ch3_x0y1,
                aib11_ch3_x0y1, aib10_ch3_x0y1, aib9_ch3_x0y1,aib8_ch3_x0y1,
                aib7_ch3_x0y1, aib6_ch3_x0y1, aib5_ch3_x0y1,aib4_ch3_x0y1,
                aib3_ch3_x0y1, aib2_ch3_x0y1, aib1_ch3_x0y1,aib0_ch3_x0y1;
    wire        aib95_ch4_x0y1, aib94_ch4_x0y1, aib93_ch4_x0y1,aib92_ch4_x0y1,
                aib91_ch4_x0y1, aib90_ch4_x0y1, aib89_ch4_x0y1,aib88_ch4_x0y1,
                aib87_ch4_x0y1, aib86_ch4_x0y1, aib85_ch4_x0y1,aib84_ch4_x0y1,
                aib83_ch4_x0y1, aib82_ch4_x0y1, aib81_ch4_x0y1,aib80_ch4_x0y1,
                aib79_ch4_x0y1, aib78_ch4_x0y1, aib77_ch4_x0y1,aib76_ch4_x0y1,
                aib75_ch4_x0y1, aib74_ch4_x0y1, aib73_ch4_x0y1,aib72_ch4_x0y1,
                aib71_ch4_x0y1, aib70_ch4_x0y1, aib69_ch4_x0y1,aib68_ch4_x0y1,
                aib67_ch4_x0y1, aib66_ch4_x0y1, aib65_ch4_x0y1,aib64_ch4_x0y1,
                aib63_ch4_x0y1, aib62_ch4_x0y1, aib61_ch4_x0y1,aib60_ch4_x0y1,
                aib59_ch4_x0y1, aib58_ch4_x0y1, aib57_ch4_x0y1,aib56_ch4_x0y1,
                aib55_ch4_x0y1, aib54_ch4_x0y1, aib53_ch4_x0y1,aib52_ch4_x0y1,
                aib51_ch4_x0y1, aib50_ch4_x0y1, aib49_ch4_x0y1,aib48_ch4_x0y1,
                aib47_ch4_x0y1, aib46_ch4_x0y1, aib45_ch4_x0y1,aib44_ch4_x0y1,
                aib43_ch4_x0y1, aib42_ch4_x0y1, aib41_ch4_x0y1,aib40_ch4_x0y1,
                aib39_ch4_x0y1, aib38_ch4_x0y1, aib37_ch4_x0y1,aib36_ch4_x0y1,
                aib35_ch4_x0y1, aib34_ch4_x0y1, aib33_ch4_x0y1,aib32_ch4_x0y1,
                aib31_ch4_x0y1, aib30_ch4_x0y1, aib29_ch4_x0y1,aib28_ch4_x0y1,
                aib27_ch4_x0y1, aib26_ch4_x0y1, aib25_ch4_x0y1,aib24_ch4_x0y1,
                aib23_ch4_x0y1, aib22_ch4_x0y1, aib21_ch4_x0y1,aib20_ch4_x0y1,
                aib19_ch4_x0y1, aib18_ch4_x0y1, aib17_ch4_x0y1,aib16_ch4_x0y1,
                aib15_ch4_x0y1, aib14_ch4_x0y1, aib13_ch4_x0y1,aib12_ch4_x0y1,
                aib11_ch4_x0y1, aib10_ch4_x0y1, aib9_ch4_x0y1,aib8_ch4_x0y1,
                aib7_ch4_x0y1, aib6_ch4_x0y1, aib5_ch4_x0y1,aib4_ch4_x0y1,
                aib3_ch4_x0y1, aib2_ch4_x0y1, aib1_ch4_x0y1,aib0_ch4_x0y1; 
    wire        aib95_ch5_x0y1, aib94_ch5_x0y1, aib93_ch5_x0y1,aib92_ch5_x0y1,
                aib91_ch5_x0y1, aib90_ch5_x0y1, aib89_ch5_x0y1,aib88_ch5_x0y1,
                aib87_ch5_x0y1, aib86_ch5_x0y1, aib85_ch5_x0y1,aib84_ch5_x0y1,
                aib83_ch5_x0y1, aib82_ch5_x0y1, aib81_ch5_x0y1,aib80_ch5_x0y1,
                aib79_ch5_x0y1, aib78_ch5_x0y1, aib77_ch5_x0y1,aib76_ch5_x0y1,
                aib75_ch5_x0y1, aib74_ch5_x0y1, aib73_ch5_x0y1,aib72_ch5_x0y1,
                aib71_ch5_x0y1, aib70_ch5_x0y1, aib69_ch5_x0y1,aib68_ch5_x0y1,
                aib67_ch5_x0y1, aib66_ch5_x0y1, aib65_ch5_x0y1,aib64_ch5_x0y1,
                aib63_ch5_x0y1, aib62_ch5_x0y1, aib61_ch5_x0y1,aib60_ch5_x0y1,
                aib59_ch5_x0y1, aib58_ch5_x0y1, aib57_ch5_x0y1,aib56_ch5_x0y1,
                aib55_ch5_x0y1, aib54_ch5_x0y1, aib53_ch5_x0y1,aib52_ch5_x0y1,
                aib51_ch5_x0y1, aib50_ch5_x0y1, aib49_ch5_x0y1,aib48_ch5_x0y1,
                aib47_ch5_x0y1, aib46_ch5_x0y1, aib45_ch5_x0y1,aib44_ch5_x0y1,
                aib43_ch5_x0y1, aib42_ch5_x0y1, aib41_ch5_x0y1,aib40_ch5_x0y1,
                aib39_ch5_x0y1, aib38_ch5_x0y1, aib37_ch5_x0y1,aib36_ch5_x0y1,
                aib35_ch5_x0y1, aib34_ch5_x0y1, aib33_ch5_x0y1,aib32_ch5_x0y1,
                aib31_ch5_x0y1, aib30_ch5_x0y1, aib29_ch5_x0y1,aib28_ch5_x0y1,
                aib27_ch5_x0y1, aib26_ch5_x0y1, aib25_ch5_x0y1,aib24_ch5_x0y1,
                aib23_ch5_x0y1, aib22_ch5_x0y1, aib21_ch5_x0y1,aib20_ch5_x0y1,
                aib19_ch5_x0y1, aib18_ch5_x0y1, aib17_ch5_x0y1,aib16_ch5_x0y1,
                aib15_ch5_x0y1, aib14_ch5_x0y1, aib13_ch5_x0y1,aib12_ch5_x0y1,
                aib11_ch5_x0y1, aib10_ch5_x0y1, aib9_ch5_x0y1,aib8_ch5_x0y1,
                aib7_ch5_x0y1, aib6_ch5_x0y1, aib5_ch5_x0y1,aib4_ch5_x0y1,
                aib3_ch5_x0y1, aib2_ch5_x0y1, aib1_ch5_x0y1,aib0_ch5_x0y1;
    wire        aib95_ch0_x0y2, aib94_ch0_x0y2, aib93_ch0_x0y2,aib92_ch0_x0y2,
                aib91_ch0_x0y2, aib90_ch0_x0y2, aib89_ch0_x0y2,aib88_ch0_x0y2,
                aib87_ch0_x0y2, aib86_ch0_x0y2, aib85_ch0_x0y2,aib84_ch0_x0y2,
                aib83_ch0_x0y2, aib82_ch0_x0y2, aib81_ch0_x0y2,aib80_ch0_x0y2,
                aib79_ch0_x0y2, aib78_ch0_x0y2, aib77_ch0_x0y2,aib76_ch0_x0y2,
                aib75_ch0_x0y2, aib74_ch0_x0y2, aib73_ch0_x0y2,aib72_ch0_x0y2,
                aib71_ch0_x0y2, aib70_ch0_x0y2, aib69_ch0_x0y2,aib68_ch0_x0y2,
                aib67_ch0_x0y2, aib66_ch0_x0y2, aib65_ch0_x0y2,aib64_ch0_x0y2,
                aib63_ch0_x0y2, aib62_ch0_x0y2, aib61_ch0_x0y2,aib60_ch0_x0y2,
                aib59_ch0_x0y2, aib58_ch0_x0y2, aib57_ch0_x0y2,aib56_ch0_x0y2,
                aib55_ch0_x0y2, aib54_ch0_x0y2, aib53_ch0_x0y2,aib52_ch0_x0y2,
                aib51_ch0_x0y2, aib50_ch0_x0y2, aib49_ch0_x0y2,aib48_ch0_x0y2,
                aib47_ch0_x0y2, aib46_ch0_x0y2, aib45_ch0_x0y2,aib44_ch0_x0y2,
                aib43_ch0_x0y2, aib42_ch0_x0y2, aib41_ch0_x0y2,aib40_ch0_x0y2,
                aib39_ch0_x0y2, aib38_ch0_x0y2, aib37_ch0_x0y2,aib36_ch0_x0y2,
                aib35_ch0_x0y2, aib34_ch0_x0y2, aib33_ch0_x0y2,aib32_ch0_x0y2,
                aib31_ch0_x0y2, aib30_ch0_x0y2, aib29_ch0_x0y2,aib28_ch0_x0y2,
                aib27_ch0_x0y2, aib26_ch0_x0y2, aib25_ch0_x0y2,aib24_ch0_x0y2,
                aib23_ch0_x0y2, aib22_ch0_x0y2, aib21_ch0_x0y2,aib20_ch0_x0y2,
                aib19_ch0_x0y2, aib18_ch0_x0y2, aib17_ch0_x0y2,aib16_ch0_x0y2,
                aib15_ch0_x0y2, aib14_ch0_x0y2, aib13_ch0_x0y2,aib12_ch0_x0y2,
                aib11_ch0_x0y2, aib10_ch0_x0y2, aib9_ch0_x0y2,aib8_ch0_x0y2,
                aib7_ch0_x0y2, aib6_ch0_x0y2, aib5_ch0_x0y2,aib4_ch0_x0y2,
                aib3_ch0_x0y2, aib2_ch0_x0y2, aib1_ch0_x0y2,aib0_ch0_x0y2;
                
    wire        aib95_ch1_x0y2, aib94_ch1_x0y2, aib93_ch1_x0y2,aib92_ch1_x0y2,
                aib91_ch1_x0y2, aib90_ch1_x0y2, aib89_ch1_x0y2,aib88_ch1_x0y2,
                aib87_ch1_x0y2, aib86_ch1_x0y2, aib85_ch1_x0y2,aib84_ch1_x0y2,
                aib83_ch1_x0y2, aib82_ch1_x0y2, aib81_ch1_x0y2,aib80_ch1_x0y2,
                aib79_ch1_x0y2, aib78_ch1_x0y2, aib77_ch1_x0y2,aib76_ch1_x0y2,
                aib75_ch1_x0y2, aib74_ch1_x0y2, aib73_ch1_x0y2,aib72_ch1_x0y2,
                aib71_ch1_x0y2, aib70_ch1_x0y2, aib69_ch1_x0y2,aib68_ch1_x0y2,
                aib67_ch1_x0y2, aib66_ch1_x0y2, aib65_ch1_x0y2,aib64_ch1_x0y2,
                aib63_ch1_x0y2, aib62_ch1_x0y2, aib61_ch1_x0y2,aib60_ch1_x0y2,
                aib59_ch1_x0y2, aib58_ch1_x0y2, aib57_ch1_x0y2,aib56_ch1_x0y2,
                aib55_ch1_x0y2, aib54_ch1_x0y2, aib53_ch1_x0y2,aib52_ch1_x0y2,
                aib51_ch1_x0y2, aib50_ch1_x0y2, aib49_ch1_x0y2,aib48_ch1_x0y2,
                aib47_ch1_x0y2, aib46_ch1_x0y2, aib45_ch1_x0y2,aib44_ch1_x0y2,
                aib43_ch1_x0y2, aib42_ch1_x0y2, aib41_ch1_x0y2,aib40_ch1_x0y2,
                aib39_ch1_x0y2, aib38_ch1_x0y2, aib37_ch1_x0y2,aib36_ch1_x0y2,
                aib35_ch1_x0y2, aib34_ch1_x0y2, aib33_ch1_x0y2,aib32_ch1_x0y2,
                aib31_ch1_x0y2, aib30_ch1_x0y2, aib29_ch1_x0y2,aib28_ch1_x0y2,
                aib27_ch1_x0y2, aib26_ch1_x0y2, aib25_ch1_x0y2,aib24_ch1_x0y2,
                aib23_ch1_x0y2, aib22_ch1_x0y2, aib21_ch1_x0y2,aib20_ch1_x0y2,
                aib19_ch1_x0y2, aib18_ch1_x0y2, aib17_ch1_x0y2,aib16_ch1_x0y2,
                aib15_ch1_x0y2, aib14_ch1_x0y2, aib13_ch1_x0y2,aib12_ch1_x0y2,
                aib11_ch1_x0y2, aib10_ch1_x0y2, aib9_ch1_x0y2,aib8_ch1_x0y2,
                aib7_ch1_x0y2, aib6_ch1_x0y2, aib5_ch1_x0y2,aib4_ch1_x0y2,
                aib3_ch1_x0y2, aib2_ch1_x0y2, aib1_ch1_x0y2,aib0_ch1_x0y2;
    wire        aib95_ch2_x0y2, aib94_ch2_x0y2, aib93_ch2_x0y2,aib92_ch2_x0y2,
                aib91_ch2_x0y2, aib90_ch2_x0y2, aib89_ch2_x0y2,aib88_ch2_x0y2,
                aib87_ch2_x0y2, aib86_ch2_x0y2, aib85_ch2_x0y2,aib84_ch2_x0y2,
                aib83_ch2_x0y2, aib82_ch2_x0y2, aib81_ch2_x0y2,aib80_ch2_x0y2,
                aib79_ch2_x0y2, aib78_ch2_x0y2, aib77_ch2_x0y2,aib76_ch2_x0y2,
                aib75_ch2_x0y2, aib74_ch2_x0y2, aib73_ch2_x0y2,aib72_ch2_x0y2,
                aib71_ch2_x0y2, aib70_ch2_x0y2, aib69_ch2_x0y2,aib68_ch2_x0y2,
                aib67_ch2_x0y2, aib66_ch2_x0y2, aib65_ch2_x0y2,aib64_ch2_x0y2,
                aib63_ch2_x0y2, aib62_ch2_x0y2, aib61_ch2_x0y2,aib60_ch2_x0y2,
                aib59_ch2_x0y2, aib58_ch2_x0y2, aib57_ch2_x0y2,aib56_ch2_x0y2,
                aib55_ch2_x0y2, aib54_ch2_x0y2, aib53_ch2_x0y2,aib52_ch2_x0y2,
                aib51_ch2_x0y2, aib50_ch2_x0y2, aib49_ch2_x0y2,aib48_ch2_x0y2,
                aib47_ch2_x0y2, aib46_ch2_x0y2, aib45_ch2_x0y2,aib44_ch2_x0y2,
                aib43_ch2_x0y2, aib42_ch2_x0y2, aib41_ch2_x0y2,aib40_ch2_x0y2,
                aib39_ch2_x0y2, aib38_ch2_x0y2, aib37_ch2_x0y2,aib36_ch2_x0y2,
                aib35_ch2_x0y2, aib34_ch2_x0y2, aib33_ch2_x0y2,aib32_ch2_x0y2,
                aib31_ch2_x0y2, aib30_ch2_x0y2, aib29_ch2_x0y2,aib28_ch2_x0y2,
                aib27_ch2_x0y2, aib26_ch2_x0y2, aib25_ch2_x0y2,aib24_ch2_x0y2,
                aib23_ch2_x0y2, aib22_ch2_x0y2, aib21_ch2_x0y2,aib20_ch2_x0y2,
                aib19_ch2_x0y2, aib18_ch2_x0y2, aib17_ch2_x0y2,aib16_ch2_x0y2,
                aib15_ch2_x0y2, aib14_ch2_x0y2, aib13_ch2_x0y2,aib12_ch2_x0y2,
                aib11_ch2_x0y2, aib10_ch2_x0y2, aib9_ch2_x0y2,aib8_ch2_x0y2,
                aib7_ch2_x0y2, aib6_ch2_x0y2, aib5_ch2_x0y2,aib4_ch2_x0y2,
                aib3_ch2_x0y2, aib2_ch2_x0y2, aib1_ch2_x0y2,aib0_ch2_x0y2; 
    wire        aib95_ch3_x0y2, aib94_ch3_x0y2, aib93_ch3_x0y2,aib92_ch3_x0y2,
                aib91_ch3_x0y2, aib90_ch3_x0y2, aib89_ch3_x0y2,aib88_ch3_x0y2,
                aib87_ch3_x0y2, aib86_ch3_x0y2, aib85_ch3_x0y2,aib84_ch3_x0y2,
                aib83_ch3_x0y2, aib82_ch3_x0y2, aib81_ch3_x0y2,aib80_ch3_x0y2,
                aib79_ch3_x0y2, aib78_ch3_x0y2, aib77_ch3_x0y2,aib76_ch3_x0y2,
                aib75_ch3_x0y2, aib74_ch3_x0y2, aib73_ch3_x0y2,aib72_ch3_x0y2,
                aib71_ch3_x0y2, aib70_ch3_x0y2, aib69_ch3_x0y2,aib68_ch3_x0y2,
                aib67_ch3_x0y2, aib66_ch3_x0y2, aib65_ch3_x0y2,aib64_ch3_x0y2,
                aib63_ch3_x0y2, aib62_ch3_x0y2, aib61_ch3_x0y2,aib60_ch3_x0y2,
                aib59_ch3_x0y2, aib58_ch3_x0y2, aib57_ch3_x0y2,aib56_ch3_x0y2,
                aib55_ch3_x0y2, aib54_ch3_x0y2, aib53_ch3_x0y2,aib52_ch3_x0y2,
                aib51_ch3_x0y2, aib50_ch3_x0y2, aib49_ch3_x0y2,aib48_ch3_x0y2,
                aib47_ch3_x0y2, aib46_ch3_x0y2, aib45_ch3_x0y2,aib44_ch3_x0y2,
                aib43_ch3_x0y2, aib42_ch3_x0y2, aib41_ch3_x0y2,aib40_ch3_x0y2,
                aib39_ch3_x0y2, aib38_ch3_x0y2, aib37_ch3_x0y2,aib36_ch3_x0y2,
                aib35_ch3_x0y2, aib34_ch3_x0y2, aib33_ch3_x0y2,aib32_ch3_x0y2,
                aib31_ch3_x0y2, aib30_ch3_x0y2, aib29_ch3_x0y2,aib28_ch3_x0y2,
                aib27_ch3_x0y2, aib26_ch3_x0y2, aib25_ch3_x0y2,aib24_ch3_x0y2,
                aib23_ch3_x0y2, aib22_ch3_x0y2, aib21_ch3_x0y2,aib20_ch3_x0y2,
                aib19_ch3_x0y2, aib18_ch3_x0y2, aib17_ch3_x0y2,aib16_ch3_x0y2,
                aib15_ch3_x0y2, aib14_ch3_x0y2, aib13_ch3_x0y2,aib12_ch3_x0y2,
                aib11_ch3_x0y2, aib10_ch3_x0y2, aib9_ch3_x0y2,aib8_ch3_x0y2,
                aib7_ch3_x0y2, aib6_ch3_x0y2, aib5_ch3_x0y2,aib4_ch3_x0y2,
                aib3_ch3_x0y2, aib2_ch3_x0y2, aib1_ch3_x0y2,aib0_ch3_x0y2;
    wire        aib95_ch4_x0y2, aib94_ch4_x0y2, aib93_ch4_x0y2,aib92_ch4_x0y2,
                aib91_ch4_x0y2, aib90_ch4_x0y2, aib89_ch4_x0y2,aib88_ch4_x0y2,
                aib87_ch4_x0y2, aib86_ch4_x0y2, aib85_ch4_x0y2,aib84_ch4_x0y2,
                aib83_ch4_x0y2, aib82_ch4_x0y2, aib81_ch4_x0y2,aib80_ch4_x0y2,
                aib79_ch4_x0y2, aib78_ch4_x0y2, aib77_ch4_x0y2,aib76_ch4_x0y2,
                aib75_ch4_x0y2, aib74_ch4_x0y2, aib73_ch4_x0y2,aib72_ch4_x0y2,
                aib71_ch4_x0y2, aib70_ch4_x0y2, aib69_ch4_x0y2,aib68_ch4_x0y2,
                aib67_ch4_x0y2, aib66_ch4_x0y2, aib65_ch4_x0y2,aib64_ch4_x0y2,
                aib63_ch4_x0y2, aib62_ch4_x0y2, aib61_ch4_x0y2,aib60_ch4_x0y2,
                aib59_ch4_x0y2, aib58_ch4_x0y2, aib57_ch4_x0y2,aib56_ch4_x0y2,
                aib55_ch4_x0y2, aib54_ch4_x0y2, aib53_ch4_x0y2,aib52_ch4_x0y2,
                aib51_ch4_x0y2, aib50_ch4_x0y2, aib49_ch4_x0y2,aib48_ch4_x0y2,
                aib47_ch4_x0y2, aib46_ch4_x0y2, aib45_ch4_x0y2,aib44_ch4_x0y2,
                aib43_ch4_x0y2, aib42_ch4_x0y2, aib41_ch4_x0y2,aib40_ch4_x0y2,
                aib39_ch4_x0y2, aib38_ch4_x0y2, aib37_ch4_x0y2,aib36_ch4_x0y2,
                aib35_ch4_x0y2, aib34_ch4_x0y2, aib33_ch4_x0y2,aib32_ch4_x0y2,
                aib31_ch4_x0y2, aib30_ch4_x0y2, aib29_ch4_x0y2,aib28_ch4_x0y2,
                aib27_ch4_x0y2, aib26_ch4_x0y2, aib25_ch4_x0y2,aib24_ch4_x0y2,
                aib23_ch4_x0y2, aib22_ch4_x0y2, aib21_ch4_x0y2,aib20_ch4_x0y2,
                aib19_ch4_x0y2, aib18_ch4_x0y2, aib17_ch4_x0y2,aib16_ch4_x0y2,
                aib15_ch4_x0y2, aib14_ch4_x0y2, aib13_ch4_x0y2,aib12_ch4_x0y2,
                aib11_ch4_x0y2, aib10_ch4_x0y2, aib9_ch4_x0y2,aib8_ch4_x0y2,
                aib7_ch4_x0y2, aib6_ch4_x0y2, aib5_ch4_x0y2,aib4_ch4_x0y2,
                aib3_ch4_x0y2, aib2_ch4_x0y2, aib1_ch4_x0y2,aib0_ch4_x0y2; 
    wire        aib95_ch5_x0y2, aib94_ch5_x0y2, aib93_ch5_x0y2,aib92_ch5_x0y2,
                aib91_ch5_x0y2, aib90_ch5_x0y2, aib89_ch5_x0y2,aib88_ch5_x0y2,
                aib87_ch5_x0y2, aib86_ch5_x0y2, aib85_ch5_x0y2,aib84_ch5_x0y2,
                aib83_ch5_x0y2, aib82_ch5_x0y2, aib81_ch5_x0y2,aib80_ch5_x0y2,
                aib79_ch5_x0y2, aib78_ch5_x0y2, aib77_ch5_x0y2,aib76_ch5_x0y2,
                aib75_ch5_x0y2, aib74_ch5_x0y2, aib73_ch5_x0y2,aib72_ch5_x0y2,
                aib71_ch5_x0y2, aib70_ch5_x0y2, aib69_ch5_x0y2,aib68_ch5_x0y2,
                aib67_ch5_x0y2, aib66_ch5_x0y2, aib65_ch5_x0y2,aib64_ch5_x0y2,
                aib63_ch5_x0y2, aib62_ch5_x0y2, aib61_ch5_x0y2,aib60_ch5_x0y2,
                aib59_ch5_x0y2, aib58_ch5_x0y2, aib57_ch5_x0y2,aib56_ch5_x0y2,
                aib55_ch5_x0y2, aib54_ch5_x0y2, aib53_ch5_x0y2,aib52_ch5_x0y2,
                aib51_ch5_x0y2, aib50_ch5_x0y2, aib49_ch5_x0y2,aib48_ch5_x0y2,
                aib47_ch5_x0y2, aib46_ch5_x0y2, aib45_ch5_x0y2,aib44_ch5_x0y2,
                aib43_ch5_x0y2, aib42_ch5_x0y2, aib41_ch5_x0y2,aib40_ch5_x0y2,
                aib39_ch5_x0y2, aib38_ch5_x0y2, aib37_ch5_x0y2,aib36_ch5_x0y2,
                aib35_ch5_x0y2, aib34_ch5_x0y2, aib33_ch5_x0y2,aib32_ch5_x0y2,
                aib31_ch5_x0y2, aib30_ch5_x0y2, aib29_ch5_x0y2,aib28_ch5_x0y2,
                aib27_ch5_x0y2, aib26_ch5_x0y2, aib25_ch5_x0y2,aib24_ch5_x0y2,
                aib23_ch5_x0y2, aib22_ch5_x0y2, aib21_ch5_x0y2,aib20_ch5_x0y2,
                aib19_ch5_x0y2, aib18_ch5_x0y2, aib17_ch5_x0y2,aib16_ch5_x0y2,
                aib15_ch5_x0y2, aib14_ch5_x0y2, aib13_ch5_x0y2,aib12_ch5_x0y2,
                aib11_ch5_x0y2, aib10_ch5_x0y2, aib9_ch5_x0y2,aib8_ch5_x0y2,
                aib7_ch5_x0y2, aib6_ch5_x0y2, aib5_ch5_x0y2,aib4_ch5_x0y2,
                aib3_ch5_x0y2, aib2_ch5_x0y2, aib1_ch5_x0y2,aib0_ch5_x0y2;
    wire        aib95_ch0_x0y3, aib94_ch0_x0y3, aib93_ch0_x0y3,aib92_ch0_x0y3,
                aib91_ch0_x0y3, aib90_ch0_x0y3, aib89_ch0_x0y3,aib88_ch0_x0y3,
                aib87_ch0_x0y3, aib86_ch0_x0y3, aib85_ch0_x0y3,aib84_ch0_x0y3,
                aib83_ch0_x0y3, aib82_ch0_x0y3, aib81_ch0_x0y3,aib80_ch0_x0y3,
                aib79_ch0_x0y3, aib78_ch0_x0y3, aib77_ch0_x0y3,aib76_ch0_x0y3,
                aib75_ch0_x0y3, aib74_ch0_x0y3, aib73_ch0_x0y3,aib72_ch0_x0y3,
                aib71_ch0_x0y3, aib70_ch0_x0y3, aib69_ch0_x0y3,aib68_ch0_x0y3,
                aib67_ch0_x0y3, aib66_ch0_x0y3, aib65_ch0_x0y3,aib64_ch0_x0y3,
                aib63_ch0_x0y3, aib62_ch0_x0y3, aib61_ch0_x0y3,aib60_ch0_x0y3,
                aib59_ch0_x0y3, aib58_ch0_x0y3, aib57_ch0_x0y3,aib56_ch0_x0y3,
                aib55_ch0_x0y3, aib54_ch0_x0y3, aib53_ch0_x0y3,aib52_ch0_x0y3,
                aib51_ch0_x0y3, aib50_ch0_x0y3, aib49_ch0_x0y3,aib48_ch0_x0y3,
                aib47_ch0_x0y3, aib46_ch0_x0y3, aib45_ch0_x0y3,aib44_ch0_x0y3,
                aib43_ch0_x0y3, aib42_ch0_x0y3, aib41_ch0_x0y3,aib40_ch0_x0y3,
                aib39_ch0_x0y3, aib38_ch0_x0y3, aib37_ch0_x0y3,aib36_ch0_x0y3,
                aib35_ch0_x0y3, aib34_ch0_x0y3, aib33_ch0_x0y3,aib32_ch0_x0y3,
                aib31_ch0_x0y3, aib30_ch0_x0y3, aib29_ch0_x0y3,aib28_ch0_x0y3,
                aib27_ch0_x0y3, aib26_ch0_x0y3, aib25_ch0_x0y3,aib24_ch0_x0y3,
                aib23_ch0_x0y3, aib22_ch0_x0y3, aib21_ch0_x0y3,aib20_ch0_x0y3,
                aib19_ch0_x0y3, aib18_ch0_x0y3, aib17_ch0_x0y3,aib16_ch0_x0y3,
                aib15_ch0_x0y3, aib14_ch0_x0y3, aib13_ch0_x0y3,aib12_ch0_x0y3,
                aib11_ch0_x0y3, aib10_ch0_x0y3, aib9_ch0_x0y3,aib8_ch0_x0y3,
                aib7_ch0_x0y3, aib6_ch0_x0y3, aib5_ch0_x0y3,aib4_ch0_x0y3,
                aib3_ch0_x0y3, aib2_ch0_x0y3, aib1_ch0_x0y3,aib0_ch0_x0y3;
                
    wire        aib95_ch1_x0y3, aib94_ch1_x0y3, aib93_ch1_x0y3,aib92_ch1_x0y3,
                aib91_ch1_x0y3, aib90_ch1_x0y3, aib89_ch1_x0y3,aib88_ch1_x0y3,
                aib87_ch1_x0y3, aib86_ch1_x0y3, aib85_ch1_x0y3,aib84_ch1_x0y3,
                aib83_ch1_x0y3, aib82_ch1_x0y3, aib81_ch1_x0y3,aib80_ch1_x0y3,
                aib79_ch1_x0y3, aib78_ch1_x0y3, aib77_ch1_x0y3,aib76_ch1_x0y3,
                aib75_ch1_x0y3, aib74_ch1_x0y3, aib73_ch1_x0y3,aib72_ch1_x0y3,
                aib71_ch1_x0y3, aib70_ch1_x0y3, aib69_ch1_x0y3,aib68_ch1_x0y3,
                aib67_ch1_x0y3, aib66_ch1_x0y3, aib65_ch1_x0y3,aib64_ch1_x0y3,
                aib63_ch1_x0y3, aib62_ch1_x0y3, aib61_ch1_x0y3,aib60_ch1_x0y3,
                aib59_ch1_x0y3, aib58_ch1_x0y3, aib57_ch1_x0y3,aib56_ch1_x0y3,
                aib55_ch1_x0y3, aib54_ch1_x0y3, aib53_ch1_x0y3,aib52_ch1_x0y3,
                aib51_ch1_x0y3, aib50_ch1_x0y3, aib49_ch1_x0y3,aib48_ch1_x0y3,
                aib47_ch1_x0y3, aib46_ch1_x0y3, aib45_ch1_x0y3,aib44_ch1_x0y3,
                aib43_ch1_x0y3, aib42_ch1_x0y3, aib41_ch1_x0y3,aib40_ch1_x0y3,
                aib39_ch1_x0y3, aib38_ch1_x0y3, aib37_ch1_x0y3,aib36_ch1_x0y3,
                aib35_ch1_x0y3, aib34_ch1_x0y3, aib33_ch1_x0y3,aib32_ch1_x0y3,
                aib31_ch1_x0y3, aib30_ch1_x0y3, aib29_ch1_x0y3,aib28_ch1_x0y3,
                aib27_ch1_x0y3, aib26_ch1_x0y3, aib25_ch1_x0y3,aib24_ch1_x0y3,
                aib23_ch1_x0y3, aib22_ch1_x0y3, aib21_ch1_x0y3,aib20_ch1_x0y3,
                aib19_ch1_x0y3, aib18_ch1_x0y3, aib17_ch1_x0y3,aib16_ch1_x0y3,
                aib15_ch1_x0y3, aib14_ch1_x0y3, aib13_ch1_x0y3,aib12_ch1_x0y3,
                aib11_ch1_x0y3, aib10_ch1_x0y3, aib9_ch1_x0y3,aib8_ch1_x0y3,
                aib7_ch1_x0y3, aib6_ch1_x0y3, aib5_ch1_x0y3,aib4_ch1_x0y3,
                aib3_ch1_x0y3, aib2_ch1_x0y3, aib1_ch1_x0y3,aib0_ch1_x0y3;
    wire        aib95_ch2_x0y3, aib94_ch2_x0y3, aib93_ch2_x0y3,aib92_ch2_x0y3,
                aib91_ch2_x0y3, aib90_ch2_x0y3, aib89_ch2_x0y3,aib88_ch2_x0y3,
                aib87_ch2_x0y3, aib86_ch2_x0y3, aib85_ch2_x0y3,aib84_ch2_x0y3,
                aib83_ch2_x0y3, aib82_ch2_x0y3, aib81_ch2_x0y3,aib80_ch2_x0y3,
                aib79_ch2_x0y3, aib78_ch2_x0y3, aib77_ch2_x0y3,aib76_ch2_x0y3,
                aib75_ch2_x0y3, aib74_ch2_x0y3, aib73_ch2_x0y3,aib72_ch2_x0y3,
                aib71_ch2_x0y3, aib70_ch2_x0y3, aib69_ch2_x0y3,aib68_ch2_x0y3,
                aib67_ch2_x0y3, aib66_ch2_x0y3, aib65_ch2_x0y3,aib64_ch2_x0y3,
                aib63_ch2_x0y3, aib62_ch2_x0y3, aib61_ch2_x0y3,aib60_ch2_x0y3,
                aib59_ch2_x0y3, aib58_ch2_x0y3, aib57_ch2_x0y3,aib56_ch2_x0y3,
                aib55_ch2_x0y3, aib54_ch2_x0y3, aib53_ch2_x0y3,aib52_ch2_x0y3,
                aib51_ch2_x0y3, aib50_ch2_x0y3, aib49_ch2_x0y3,aib48_ch2_x0y3,
                aib47_ch2_x0y3, aib46_ch2_x0y3, aib45_ch2_x0y3,aib44_ch2_x0y3,
                aib43_ch2_x0y3, aib42_ch2_x0y3, aib41_ch2_x0y3,aib40_ch2_x0y3,
                aib39_ch2_x0y3, aib38_ch2_x0y3, aib37_ch2_x0y3,aib36_ch2_x0y3,
                aib35_ch2_x0y3, aib34_ch2_x0y3, aib33_ch2_x0y3,aib32_ch2_x0y3,
                aib31_ch2_x0y3, aib30_ch2_x0y3, aib29_ch2_x0y3,aib28_ch2_x0y3,
                aib27_ch2_x0y3, aib26_ch2_x0y3, aib25_ch2_x0y3,aib24_ch2_x0y3,
                aib23_ch2_x0y3, aib22_ch2_x0y3, aib21_ch2_x0y3,aib20_ch2_x0y3,
                aib19_ch2_x0y3, aib18_ch2_x0y3, aib17_ch2_x0y3,aib16_ch2_x0y3,
                aib15_ch2_x0y3, aib14_ch2_x0y3, aib13_ch2_x0y3,aib12_ch2_x0y3,
                aib11_ch2_x0y3, aib10_ch2_x0y3, aib9_ch2_x0y3,aib8_ch2_x0y3,
                aib7_ch2_x0y3, aib6_ch2_x0y3, aib5_ch2_x0y3,aib4_ch2_x0y3,
                aib3_ch2_x0y3, aib2_ch2_x0y3, aib1_ch2_x0y3,aib0_ch2_x0y3; 
    wire        aib95_ch3_x0y3, aib94_ch3_x0y3, aib93_ch3_x0y3,aib92_ch3_x0y3,
                aib91_ch3_x0y3, aib90_ch3_x0y3, aib89_ch3_x0y3,aib88_ch3_x0y3,
                aib87_ch3_x0y3, aib86_ch3_x0y3, aib85_ch3_x0y3,aib84_ch3_x0y3,
                aib83_ch3_x0y3, aib82_ch3_x0y3, aib81_ch3_x0y3,aib80_ch3_x0y3,
                aib79_ch3_x0y3, aib78_ch3_x0y3, aib77_ch3_x0y3,aib76_ch3_x0y3,
                aib75_ch3_x0y3, aib74_ch3_x0y3, aib73_ch3_x0y3,aib72_ch3_x0y3,
                aib71_ch3_x0y3, aib70_ch3_x0y3, aib69_ch3_x0y3,aib68_ch3_x0y3,
                aib67_ch3_x0y3, aib66_ch3_x0y3, aib65_ch3_x0y3,aib64_ch3_x0y3,
                aib63_ch3_x0y3, aib62_ch3_x0y3, aib61_ch3_x0y3,aib60_ch3_x0y3,
                aib59_ch3_x0y3, aib58_ch3_x0y3, aib57_ch3_x0y3,aib56_ch3_x0y3,
                aib55_ch3_x0y3, aib54_ch3_x0y3, aib53_ch3_x0y3,aib52_ch3_x0y3,
                aib51_ch3_x0y3, aib50_ch3_x0y3, aib49_ch3_x0y3,aib48_ch3_x0y3,
                aib47_ch3_x0y3, aib46_ch3_x0y3, aib45_ch3_x0y3,aib44_ch3_x0y3,
                aib43_ch3_x0y3, aib42_ch3_x0y3, aib41_ch3_x0y3,aib40_ch3_x0y3,
                aib39_ch3_x0y3, aib38_ch3_x0y3, aib37_ch3_x0y3,aib36_ch3_x0y3,
                aib35_ch3_x0y3, aib34_ch3_x0y3, aib33_ch3_x0y3,aib32_ch3_x0y3,
                aib31_ch3_x0y3, aib30_ch3_x0y3, aib29_ch3_x0y3,aib28_ch3_x0y3,
                aib27_ch3_x0y3, aib26_ch3_x0y3, aib25_ch3_x0y3,aib24_ch3_x0y3,
                aib23_ch3_x0y3, aib22_ch3_x0y3, aib21_ch3_x0y3,aib20_ch3_x0y3,
                aib19_ch3_x0y3, aib18_ch3_x0y3, aib17_ch3_x0y3,aib16_ch3_x0y3,
                aib15_ch3_x0y3, aib14_ch3_x0y3, aib13_ch3_x0y3,aib12_ch3_x0y3,
                aib11_ch3_x0y3, aib10_ch3_x0y3, aib9_ch3_x0y3,aib8_ch3_x0y3,
                aib7_ch3_x0y3, aib6_ch3_x0y3, aib5_ch3_x0y3,aib4_ch3_x0y3,
                aib3_ch3_x0y3, aib2_ch3_x0y3, aib1_ch3_x0y3,aib0_ch3_x0y3;
    wire        aib95_ch4_x0y3, aib94_ch4_x0y3, aib93_ch4_x0y3,aib92_ch4_x0y3,
                aib91_ch4_x0y3, aib90_ch4_x0y3, aib89_ch4_x0y3,aib88_ch4_x0y3,
                aib87_ch4_x0y3, aib86_ch4_x0y3, aib85_ch4_x0y3,aib84_ch4_x0y3,
                aib83_ch4_x0y3, aib82_ch4_x0y3, aib81_ch4_x0y3,aib80_ch4_x0y3,
                aib79_ch4_x0y3, aib78_ch4_x0y3, aib77_ch4_x0y3,aib76_ch4_x0y3,
                aib75_ch4_x0y3, aib74_ch4_x0y3, aib73_ch4_x0y3,aib72_ch4_x0y3,
                aib71_ch4_x0y3, aib70_ch4_x0y3, aib69_ch4_x0y3,aib68_ch4_x0y3,
                aib67_ch4_x0y3, aib66_ch4_x0y3, aib65_ch4_x0y3,aib64_ch4_x0y3,
                aib63_ch4_x0y3, aib62_ch4_x0y3, aib61_ch4_x0y3,aib60_ch4_x0y3,
                aib59_ch4_x0y3, aib58_ch4_x0y3, aib57_ch4_x0y3,aib56_ch4_x0y3,
                aib55_ch4_x0y3, aib54_ch4_x0y3, aib53_ch4_x0y3,aib52_ch4_x0y3,
                aib51_ch4_x0y3, aib50_ch4_x0y3, aib49_ch4_x0y3,aib48_ch4_x0y3,
                aib47_ch4_x0y3, aib46_ch4_x0y3, aib45_ch4_x0y3,aib44_ch4_x0y3,
                aib43_ch4_x0y3, aib42_ch4_x0y3, aib41_ch4_x0y3,aib40_ch4_x0y3,
                aib39_ch4_x0y3, aib38_ch4_x0y3, aib37_ch4_x0y3,aib36_ch4_x0y3,
                aib35_ch4_x0y3, aib34_ch4_x0y3, aib33_ch4_x0y3,aib32_ch4_x0y3,
                aib31_ch4_x0y3, aib30_ch4_x0y3, aib29_ch4_x0y3,aib28_ch4_x0y3,
                aib27_ch4_x0y3, aib26_ch4_x0y3, aib25_ch4_x0y3,aib24_ch4_x0y3,
                aib23_ch4_x0y3, aib22_ch4_x0y3, aib21_ch4_x0y3,aib20_ch4_x0y3,
                aib19_ch4_x0y3, aib18_ch4_x0y3, aib17_ch4_x0y3,aib16_ch4_x0y3,
                aib15_ch4_x0y3, aib14_ch4_x0y3, aib13_ch4_x0y3,aib12_ch4_x0y3,
                aib11_ch4_x0y3, aib10_ch4_x0y3, aib9_ch4_x0y3,aib8_ch4_x0y3,
                aib7_ch4_x0y3, aib6_ch4_x0y3, aib5_ch4_x0y3,aib4_ch4_x0y3,
                aib3_ch4_x0y3, aib2_ch4_x0y3, aib1_ch4_x0y3,aib0_ch4_x0y3; 
    wire        aib95_ch5_x0y3, aib94_ch5_x0y3, aib93_ch5_x0y3,aib92_ch5_x0y3,
                aib91_ch5_x0y3, aib90_ch5_x0y3, aib89_ch5_x0y3,aib88_ch5_x0y3,
                aib87_ch5_x0y3, aib86_ch5_x0y3, aib85_ch5_x0y3,aib84_ch5_x0y3,
                aib83_ch5_x0y3, aib82_ch5_x0y3, aib81_ch5_x0y3,aib80_ch5_x0y3,
                aib79_ch5_x0y3, aib78_ch5_x0y3, aib77_ch5_x0y3,aib76_ch5_x0y3,
                aib75_ch5_x0y3, aib74_ch5_x0y3, aib73_ch5_x0y3,aib72_ch5_x0y3,
                aib71_ch5_x0y3, aib70_ch5_x0y3, aib69_ch5_x0y3,aib68_ch5_x0y3,
                aib67_ch5_x0y3, aib66_ch5_x0y3, aib65_ch5_x0y3,aib64_ch5_x0y3,
                aib63_ch5_x0y3, aib62_ch5_x0y3, aib61_ch5_x0y3,aib60_ch5_x0y3,
                aib59_ch5_x0y3, aib58_ch5_x0y3, aib57_ch5_x0y3,aib56_ch5_x0y3,
                aib55_ch5_x0y3, aib54_ch5_x0y3, aib53_ch5_x0y3,aib52_ch5_x0y3,
                aib51_ch5_x0y3, aib50_ch5_x0y3, aib49_ch5_x0y3,aib48_ch5_x0y3,
                aib47_ch5_x0y3, aib46_ch5_x0y3, aib45_ch5_x0y3,aib44_ch5_x0y3,
                aib43_ch5_x0y3, aib42_ch5_x0y3, aib41_ch5_x0y3,aib40_ch5_x0y3,
                aib39_ch5_x0y3, aib38_ch5_x0y3, aib37_ch5_x0y3,aib36_ch5_x0y3,
                aib35_ch5_x0y3, aib34_ch5_x0y3, aib33_ch5_x0y3,aib32_ch5_x0y3,
                aib31_ch5_x0y3, aib30_ch5_x0y3, aib29_ch5_x0y3,aib28_ch5_x0y3,
                aib27_ch5_x0y3, aib26_ch5_x0y3, aib25_ch5_x0y3,aib24_ch5_x0y3,
                aib23_ch5_x0y3, aib22_ch5_x0y3, aib21_ch5_x0y3,aib20_ch5_x0y3,
                aib19_ch5_x0y3, aib18_ch5_x0y3, aib17_ch5_x0y3,aib16_ch5_x0y3,
                aib15_ch5_x0y3, aib14_ch5_x0y3, aib13_ch5_x0y3,aib12_ch5_x0y3,
                aib11_ch5_x0y3, aib10_ch5_x0y3, aib9_ch5_x0y3,aib8_ch5_x0y3,
                aib7_ch5_x0y3, aib6_ch5_x0y3, aib5_ch5_x0y3,aib4_ch5_x0y3,
                aib3_ch5_x0y3, aib2_ch5_x0y3, aib1_ch5_x0y3,aib0_ch5_x0y3;
    wire        aib_aux95_x0y0, aib_aux94_x0y0, aib_aux93_x0y0,aib_aux92_x0y0,
                aib_aux91_x0y0, aib_aux90_x0y0, aib_aux89_x0y0,aib_aux88_x0y0,
                aib_aux87_x0y0, aib_aux86_x0y0, aib_aux85_x0y0,aib_aux84_x0y0,
                aib_aux83_x0y0, aib_aux82_x0y0, aib_aux81_x0y0,aib_aux80_x0y0,
                aib_aux79_x0y0, aib_aux78_x0y0, aib_aux77_x0y0,aib_aux76_x0y0,
                aib_aux75_x0y0, aib_aux74_x0y0, aib_aux73_x0y0,aib_aux72_x0y0,
                aib_aux71_x0y0, aib_aux70_x0y0, aib_aux69_x0y0,aib_aux68_x0y0,
                aib_aux67_x0y0, aib_aux66_x0y0, aib_aux65_x0y0,aib_aux64_x0y0,
                aib_aux63_x0y0, aib_aux62_x0y0, aib_aux61_x0y0,aib_aux60_x0y0,
                aib_aux59_x0y0, aib_aux58_x0y0, aib_aux57_x0y0,aib_aux56_x0y0,
                aib_aux55_x0y0, aib_aux54_x0y0, aib_aux53_x0y0,aib_aux52_x0y0,
                aib_aux51_x0y0, aib_aux50_x0y0, aib_aux49_x0y0,aib_aux48_x0y0,
                aib_aux47_x0y0, aib_aux46_x0y0, aib_aux45_x0y0,aib_aux44_x0y0,
                aib_aux43_x0y0, aib_aux42_x0y0, aib_aux41_x0y0,aib_aux40_x0y0,
                aib_aux39_x0y0, aib_aux38_x0y0, aib_aux37_x0y0,aib_aux36_x0y0,
                aib_aux35_x0y0, aib_aux34_x0y0, aib_aux33_x0y0,aib_aux32_x0y0,
                aib_aux31_x0y0, aib_aux30_x0y0, aib_aux29_x0y0,aib_aux28_x0y0,
                aib_aux27_x0y0, aib_aux26_x0y0, aib_aux25_x0y0,aib_aux24_x0y0,
                aib_aux23_x0y0, aib_aux22_x0y0, aib_aux21_x0y0,aib_aux20_x0y0,
                aib_aux19_x0y0, aib_aux18_x0y0, aib_aux17_x0y0,aib_aux16_x0y0,
                aib_aux15_x0y0, aib_aux14_x0y0, aib_aux13_x0y0,aib_aux12_x0y0,
                aib_aux11_x0y0, aib_aux10_x0y0, aib_aux9_x0y0,aib_aux8_x0y0,
                aib_aux7_x0y0, aib_aux6_x0y0, aib_aux5_x0y0,aib_aux4_x0y0,
                aib_aux3_x0y0, aib_aux2_x0y0, aib_aux1_x0y0,aib_aux0_x0y0; 
   wire [24*40-1:0] o_tx_pma_data_24ch;
// wire [39:0] o_tx_pma_data = o_tx_pma_data_24ch[39:0];

/*///////////////////////////////////////////////////////////////////////////
   aib[19:0]  loopback to aib[39:20]  --transfer data    -> receiving data
   aib[41:40] loopback to aib[43:42]  --transfer clk     -> receiving clk
   aib[85:84] loopback to aib[83:82]  --transfer sr_clk  -> receiving sr_clk
   aib[94]    loopback to aib[92]     --ssr_load_out     -> ssr_load_in

   The following pins are tied to high so that the loopback test will work:
   aib[93] -- ssr_data_in
   aib[65] -- adapter_rx_pld_rst_n
   aib[61] -- adapter_tx_pld_rst_n
   
*///////////////////////////////////////////////////////////////////////////   
/*
   assign AIB_CHAN0 = {aib95_ch0_x0y0, aib94_ch0_x0y0, 1'b1,          aib94_ch0_x0y0,
                aib91_ch0_x0y0, aib90_ch0_x0y0, aib89_ch0_x0y0,aib88_ch0_x0y0,
                aib87_ch0_x0y0, aib86_ch0_x0y0, aib85_ch0_x0y0,aib84_ch0_x0y0,
                aib85_ch0_x0y0, aib82_ch0_x0y0, aib81_ch0_x0y0,aib80_ch0_x0y0,
                aib79_ch0_x0y0, aib78_ch0_x0y0, aib77_ch0_x0y0,aib76_ch0_x0y0,
                aib75_ch0_x0y0, aib74_ch0_x0y0, aib73_ch0_x0y0,aib72_ch0_x0y0,
                aib71_ch0_x0y0, aib70_ch0_x0y0, aib69_ch0_x0y0,aib68_ch0_x0y0,
                aib67_ch0_x0y0, aib66_ch0_x0y0, 1'b1,          aib64_ch0_x0y0,
                aib63_ch0_x0y0, aib62_ch0_x0y0, 1'b1,          aib60_ch0_x0y0,
                aib59_ch0_x0y0, aib58_ch0_x0y0, aib57_ch0_x0y0,aib56_ch0_x0y0,
                aib55_ch0_x0y0, aib54_ch0_x0y0, aib53_ch0_x0y0,aib52_ch0_x0y0,
                aib51_ch0_x0y0, aib50_ch0_x0y0, aib49_ch0_x0y0,aib48_ch0_x0y0,
                aib47_ch0_x0y0, aib46_ch0_x0y0, aib45_ch0_x0y0,aib44_ch0_x0y0,
                aib41_ch0_x0y0, aib40_ch0_x0y0, aib41_ch0_x0y0,aib40_ch0_x0y0,
                aib19_ch0_x0y0, aib18_ch0_x0y0, aib17_ch0_x0y0,aib16_ch0_x0y0,
                aib15_ch0_x0y0, aib14_ch0_x0y0, aib13_ch0_x0y0,aib12_ch0_x0y0,
                aib11_ch0_x0y0, aib10_ch0_x0y0, aib9_ch0_x0y0, aib8_ch0_x0y0,
                aib7_ch0_x0y0,  aib6_ch0_x0y0,  aib5_ch0_x0y0, aib4_ch0_x0y0,
                aib3_ch0_x0y0,  aib2_ch0_x0y0,  aib1_ch0_x0y0, aib0_ch0_x0y0,
                aib19_ch0_x0y0, aib18_ch0_x0y0, aib17_ch0_x0y0,aib16_ch0_x0y0,
                aib15_ch0_x0y0, aib14_ch0_x0y0, aib13_ch0_x0y0,aib12_ch0_x0y0,
                aib11_ch0_x0y0, aib10_ch0_x0y0, aib9_ch0_x0y0, aib8_ch0_x0y0,
                aib7_ch0_x0y0,  aib6_ch0_x0y0,  aib5_ch0_x0y0, aib4_ch0_x0y0,
                aib3_ch0_x0y0,  aib2_ch0_x0y0,  aib1_ch0_x0y0, aib0_ch0_x0y0};

  assign AIB_CHAN1 = {aib95_ch1_x0y0, aib94_ch1_x0y0, 1'b1,          aib94_ch1_x0y0,
                aib91_ch1_x0y0, aib90_ch1_x0y0, aib89_ch1_x0y0,aib88_ch1_x0y0,
                aib87_ch1_x0y0, aib86_ch1_x0y0, aib85_ch1_x0y0,aib84_ch1_x0y0,
                aib85_ch1_x0y0, aib84_ch1_x0y0, aib81_ch1_x0y0,aib80_ch1_x0y0,
                aib79_ch1_x0y0, aib78_ch1_x0y0, aib77_ch1_x0y0,aib76_ch1_x0y0,
                aib75_ch1_x0y0, aib74_ch1_x0y0, aib73_ch1_x0y0,aib72_ch1_x0y0,
                aib71_ch1_x0y0, aib70_ch1_x0y0, aib69_ch1_x0y0,aib68_ch1_x0y0,
                aib67_ch1_x0y0, aib66_ch1_x0y0, 1'b1,          aib64_ch1_x0y0,
                aib63_ch1_x0y0, aib62_ch1_x0y0, 1'b1,          aib60_ch1_x0y0,
                aib59_ch1_x0y0, aib58_ch1_x0y0, aib57_ch1_x0y0,aib56_ch1_x0y0,
                aib55_ch1_x0y0, aib54_ch1_x0y0, aib53_ch1_x0y0,aib52_ch1_x0y0,
                aib51_ch1_x0y0, aib50_ch1_x0y0, aib49_ch1_x0y0,aib48_ch1_x0y0,
                aib47_ch1_x0y0, aib46_ch1_x0y0, aib45_ch1_x0y0,aib44_ch1_x0y0,
                aib41_ch1_x0y0, aib40_ch1_x0y0, aib41_ch1_x0y0,aib40_ch1_x0y0,
                aib19_ch1_x0y0, aib18_ch1_x0y0, aib17_ch1_x0y0,aib16_ch1_x0y0,
                aib15_ch1_x0y0, aib14_ch1_x0y0, aib13_ch1_x0y0,aib12_ch1_x0y0,
                aib11_ch1_x0y0, aib10_ch1_x0y0, aib9_ch1_x0y0, aib8_ch1_x0y0,
                aib7_ch1_x0y0,  aib6_ch1_x0y0,  aib5_ch1_x0y0, aib4_ch1_x0y0,
                aib3_ch1_x0y0,  aib2_ch1_x0y0,  aib1_ch1_x0y0, aib0_ch1_x0y0,
                aib19_ch1_x0y0, aib18_ch1_x0y0, aib17_ch1_x0y0,aib16_ch1_x0y0,
                aib15_ch1_x0y0, aib14_ch1_x0y0, aib13_ch1_x0y0,aib12_ch1_x0y0,
                aib11_ch1_x0y0, aib10_ch1_x0y0, aib9_ch1_x0y0, aib8_ch1_x0y0,
                aib7_ch1_x0y0,  aib6_ch1_x0y0,  aib5_ch1_x0y0, aib4_ch1_x0y0,
                aib3_ch1_x0y0,  aib2_ch1_x0y0,  aib1_ch1_x0y0, aib0_ch1_x0y0};

  assign AIB_CHAN2 = {aib95_ch2_x0y0, aib94_ch2_x0y0, 1'b1,          aib94_ch2_x0y0,
                aib91_ch2_x0y0, aib90_ch2_x0y0, aib89_ch2_x0y0,aib88_ch2_x0y0,
                aib87_ch2_x0y0, aib86_ch2_x0y0, aib85_ch2_x0y0,aib84_ch2_x0y0,
                aib85_ch2_x0y0, aib84_ch2_x0y0, aib81_ch2_x0y0,aib80_ch2_x0y0,
                aib79_ch2_x0y0, aib78_ch2_x0y0, aib77_ch2_x0y0,aib76_ch2_x0y0,
                aib75_ch2_x0y0, aib74_ch2_x0y0, aib73_ch2_x0y0,aib72_ch2_x0y0,
                aib71_ch2_x0y0, aib70_ch2_x0y0, aib69_ch2_x0y0,aib68_ch2_x0y0,
                aib67_ch2_x0y0, aib66_ch2_x0y0, 1'b1,          aib64_ch2_x0y0,
                aib63_ch2_x0y0, aib62_ch2_x0y0, 1'b1,          aib60_ch2_x0y0,
                aib59_ch2_x0y0, aib58_ch2_x0y0, aib57_ch2_x0y0,aib56_ch2_x0y0,
                aib55_ch2_x0y0, aib54_ch2_x0y0, aib53_ch2_x0y0,aib52_ch2_x0y0,
                aib51_ch2_x0y0, aib50_ch2_x0y0, aib49_ch2_x0y0,aib48_ch2_x0y0,
                aib47_ch2_x0y0, aib46_ch2_x0y0, aib45_ch2_x0y0,aib44_ch2_x0y0,
                aib41_ch2_x0y0, aib40_ch2_x0y0, aib41_ch2_x0y0,aib40_ch2_x0y0,
                aib19_ch2_x0y0, aib18_ch2_x0y0, aib17_ch2_x0y0,aib16_ch2_x0y0,
                aib15_ch2_x0y0, aib14_ch2_x0y0, aib13_ch2_x0y0,aib12_ch2_x0y0,
                aib11_ch2_x0y0, aib10_ch2_x0y0, aib9_ch2_x0y0, aib8_ch2_x0y0,
                aib7_ch2_x0y0,  aib6_ch2_x0y0,  aib5_ch2_x0y0, aib4_ch2_x0y0,
                aib3_ch2_x0y0,  aib2_ch2_x0y0,  aib1_ch2_x0y0, aib0_ch2_x0y0,
                aib19_ch2_x0y0, aib18_ch2_x0y0, aib17_ch2_x0y0,aib16_ch2_x0y0,
                aib15_ch2_x0y0, aib14_ch2_x0y0, aib13_ch2_x0y0,aib12_ch2_x0y0,
                aib11_ch2_x0y0, aib10_ch2_x0y0, aib9_ch2_x0y0, aib8_ch2_x0y0,
                aib7_ch2_x0y0,  aib6_ch2_x0y0,  aib5_ch2_x0y0, aib4_ch2_x0y0,
                aib3_ch2_x0y0,  aib2_ch2_x0y0,  aib1_ch2_x0y0, aib0_ch2_x0y0};

  assign AIB_CHAN3 = {aib95_ch3_x0y0, aib94_ch3_x0y0, 1'b1,          aib94_ch3_x0y0,
                aib91_ch3_x0y0, aib90_ch3_x0y0, aib89_ch3_x0y0,aib88_ch3_x0y0,
                aib87_ch3_x0y0, aib86_ch3_x0y0, aib85_ch3_x0y0,aib84_ch3_x0y0,
                aib85_ch3_x0y0, aib84_ch3_x0y0, aib81_ch3_x0y0,aib80_ch3_x0y0,
                aib79_ch3_x0y0, aib78_ch3_x0y0, aib77_ch3_x0y0,aib76_ch3_x0y0,
                aib75_ch3_x0y0, aib74_ch3_x0y0, aib73_ch3_x0y0,aib72_ch3_x0y0,
                aib71_ch3_x0y0, aib70_ch3_x0y0, aib69_ch3_x0y0,aib68_ch3_x0y0,
                aib67_ch3_x0y0, aib66_ch3_x0y0, 1'b1,          aib64_ch3_x0y0,
                aib63_ch3_x0y0, aib62_ch3_x0y0, 1'b1,          aib60_ch3_x0y0,
                aib59_ch3_x0y0, aib58_ch3_x0y0, aib57_ch3_x0y0,aib56_ch3_x0y0,
                aib55_ch3_x0y0, aib54_ch3_x0y0, aib53_ch3_x0y0,aib52_ch3_x0y0,
                aib51_ch3_x0y0, aib50_ch3_x0y0, aib49_ch3_x0y0,aib48_ch3_x0y0,
                aib47_ch3_x0y0, aib46_ch3_x0y0, aib45_ch3_x0y0,aib44_ch3_x0y0,
                aib41_ch3_x0y0, aib40_ch3_x0y0, aib41_ch3_x0y0,aib40_ch3_x0y0,
                aib19_ch3_x0y0, aib18_ch3_x0y0, aib17_ch3_x0y0,aib16_ch3_x0y0,
                aib15_ch3_x0y0, aib14_ch3_x0y0, aib13_ch3_x0y0,aib12_ch3_x0y0,
                aib11_ch3_x0y0, aib10_ch3_x0y0, aib9_ch3_x0y0, aib8_ch3_x0y0,
                aib7_ch3_x0y0,  aib6_ch3_x0y0,  aib5_ch3_x0y0, aib4_ch3_x0y0,
                aib3_ch3_x0y0,  aib2_ch3_x0y0,  aib1_ch3_x0y0, aib0_ch3_x0y0,
                aib19_ch3_x0y0, aib18_ch3_x0y0, aib17_ch3_x0y0,aib16_ch3_x0y0,
                aib15_ch3_x0y0, aib14_ch3_x0y0, aib13_ch3_x0y0,aib12_ch3_x0y0,
                aib11_ch3_x0y0, aib10_ch3_x0y0, aib9_ch3_x0y0, aib8_ch3_x0y0,
                aib7_ch3_x0y0,  aib6_ch3_x0y0,  aib5_ch3_x0y0, aib4_ch3_x0y0,
                aib3_ch3_x0y0,  aib2_ch3_x0y0,  aib1_ch3_x0y0, aib0_ch3_x0y0};

  assign AIB_CHAN4 = {aib95_ch4_x0y0, aib94_ch4_x0y0, 1'b1,          aib94_ch4_x0y0,
                aib91_ch4_x0y0, aib90_ch4_x0y0, aib89_ch4_x0y0,aib88_ch4_x0y0,
                aib87_ch4_x0y0, aib86_ch4_x0y0, aib85_ch4_x0y0,aib84_ch4_x0y0,
                aib85_ch4_x0y0, aib84_ch4_x0y0, aib81_ch4_x0y0,aib80_ch4_x0y0,
                aib79_ch4_x0y0, aib78_ch4_x0y0, aib77_ch4_x0y0,aib76_ch4_x0y0,
                aib75_ch4_x0y0, aib74_ch4_x0y0, aib73_ch4_x0y0,aib72_ch4_x0y0,
                aib71_ch4_x0y0, aib70_ch4_x0y0, aib69_ch4_x0y0,aib68_ch4_x0y0,
                aib67_ch4_x0y0, aib66_ch4_x0y0, 1'b1,          aib64_ch4_x0y0,
                aib63_ch4_x0y0, aib62_ch4_x0y0, 1'b1,          aib60_ch4_x0y0,
                aib59_ch4_x0y0, aib58_ch4_x0y0, aib57_ch4_x0y0,aib56_ch4_x0y0,
                aib55_ch4_x0y0, aib54_ch4_x0y0, aib53_ch4_x0y0,aib52_ch4_x0y0,
                aib51_ch4_x0y0, aib50_ch4_x0y0, aib49_ch4_x0y0,aib48_ch4_x0y0,
                aib47_ch4_x0y0, aib46_ch4_x0y0, aib45_ch4_x0y0,aib44_ch4_x0y0,
                aib41_ch4_x0y0, aib40_ch4_x0y0, aib41_ch4_x0y0,aib40_ch4_x0y0,
                aib19_ch4_x0y0, aib18_ch4_x0y0, aib17_ch4_x0y0,aib16_ch4_x0y0,
                aib15_ch4_x0y0, aib14_ch4_x0y0, aib13_ch4_x0y0,aib12_ch4_x0y0,
                aib11_ch4_x0y0, aib10_ch4_x0y0, aib9_ch4_x0y0, aib8_ch4_x0y0,
                aib7_ch4_x0y0,  aib6_ch4_x0y0,  aib5_ch4_x0y0, aib4_ch4_x0y0,
                aib3_ch4_x0y0,  aib2_ch4_x0y0,  aib1_ch4_x0y0, aib0_ch4_x0y0,
                aib19_ch4_x0y0, aib18_ch4_x0y0, aib17_ch4_x0y0,aib16_ch4_x0y0,
                aib15_ch4_x0y0, aib14_ch4_x0y0, aib13_ch4_x0y0,aib12_ch4_x0y0,
                aib11_ch4_x0y0, aib10_ch4_x0y0, aib9_ch4_x0y0, aib8_ch4_x0y0,
                aib7_ch4_x0y0,  aib6_ch4_x0y0,  aib5_ch4_x0y0, aib4_ch4_x0y0,
                aib3_ch4_x0y0,  aib2_ch4_x0y0,  aib1_ch4_x0y0, aib0_ch4_x0y0};

  assign AIB_CHAN5 = {aib95_ch5_x0y0, aib94_ch5_x0y0, 1'b1,          aib94_ch5_x0y0,
                aib91_ch5_x0y0, aib90_ch5_x0y0, aib89_ch5_x0y0,aib88_ch5_x0y0,
                aib87_ch5_x0y0, aib86_ch5_x0y0, aib85_ch5_x0y0,aib84_ch5_x0y0,
                aib85_ch5_x0y0, aib84_ch5_x0y0, aib81_ch5_x0y0,aib80_ch5_x0y0,
                aib79_ch5_x0y0, aib78_ch5_x0y0, aib77_ch5_x0y0,aib76_ch5_x0y0,
                aib75_ch5_x0y0, aib74_ch5_x0y0, aib73_ch5_x0y0,aib72_ch5_x0y0,
                aib71_ch5_x0y0, aib70_ch5_x0y0, aib69_ch5_x0y0,aib68_ch5_x0y0,
                aib67_ch5_x0y0, aib66_ch5_x0y0, 1'b1,          aib64_ch5_x0y0,
                aib63_ch5_x0y0, aib62_ch5_x0y0, 1'b1,          aib60_ch5_x0y0,
                aib59_ch5_x0y0, aib58_ch5_x0y0, aib57_ch5_x0y0,aib56_ch5_x0y0,
                aib55_ch5_x0y0, aib54_ch5_x0y0, aib53_ch5_x0y0,aib52_ch5_x0y0,
                aib51_ch5_x0y0, aib50_ch5_x0y0, aib49_ch5_x0y0,aib48_ch5_x0y0,
                aib47_ch5_x0y0, aib46_ch5_x0y0, aib45_ch5_x0y0,aib44_ch5_x0y0,
                aib41_ch5_x0y0, aib40_ch5_x0y0, aib41_ch5_x0y0,aib40_ch5_x0y0,
                aib19_ch5_x0y0, aib18_ch5_x0y0, aib17_ch5_x0y0,aib16_ch5_x0y0,
                aib15_ch5_x0y0, aib14_ch5_x0y0, aib13_ch5_x0y0,aib12_ch5_x0y0,
                aib11_ch5_x0y0, aib10_ch5_x0y0, aib9_ch5_x0y0, aib8_ch5_x0y0,
                aib7_ch5_x0y0,  aib6_ch5_x0y0,  aib5_ch5_x0y0, aib4_ch5_x0y0,
                aib3_ch5_x0y0,  aib2_ch5_x0y0,  aib1_ch5_x0y0, aib0_ch5_x0y0,
                aib19_ch5_x0y0, aib18_ch5_x0y0, aib17_ch5_x0y0,aib16_ch5_x0y0,
                aib15_ch5_x0y0, aib14_ch5_x0y0, aib13_ch5_x0y0,aib12_ch5_x0y0,
                aib11_ch5_x0y0, aib10_ch5_x0y0, aib9_ch5_x0y0, aib8_ch5_x0y0,
                aib7_ch5_x0y0,  aib6_ch5_x0y0,  aib5_ch5_x0y0, aib4_ch5_x0y0,
                aib3_ch5_x0y0,  aib2_ch5_x0y0,  aib1_ch5_x0y0, aib0_ch5_x0y0};

  assign AIB_CHAN6 = {aib95_ch0_x0y1, aib94_ch0_x0y1, 1'b1,          aib94_ch0_x0y1,
                aib91_ch0_x0y1, aib90_ch0_x0y1, aib89_ch0_x0y1,aib88_ch0_x0y1,
                aib87_ch0_x0y1, aib86_ch0_x0y1, aib85_ch0_x0y1,aib84_ch0_x0y1,
                aib85_ch0_x0y1, aib84_ch0_x0y1, aib81_ch0_x0y1,aib80_ch0_x0y1,
                aib79_ch0_x0y1, aib78_ch0_x0y1, aib77_ch0_x0y1,aib76_ch0_x0y1,
                aib75_ch0_x0y1, aib74_ch0_x0y1, aib73_ch0_x0y1,aib72_ch0_x0y1,
                aib71_ch0_x0y1, aib70_ch0_x0y1, aib69_ch0_x0y1,aib68_ch0_x0y1,
                aib67_ch0_x0y1, aib66_ch0_x0y1, 1'b1,          aib64_ch0_x0y1,
                aib63_ch0_x0y1, aib62_ch0_x0y1, 1'b1,          aib60_ch0_x0y1,
                aib59_ch0_x0y1, aib58_ch0_x0y1, aib57_ch0_x0y1,aib56_ch0_x0y1,
                aib55_ch0_x0y1, aib54_ch0_x0y1, aib53_ch0_x0y1,aib52_ch0_x0y1,
                aib51_ch0_x0y1, aib50_ch0_x0y1, aib49_ch0_x0y1,aib48_ch0_x0y1,
                aib47_ch0_x0y1, aib46_ch0_x0y1, aib45_ch0_x0y1,aib44_ch0_x0y1,
                aib41_ch0_x0y1, aib40_ch0_x0y1, aib41_ch0_x0y1,aib40_ch0_x0y1,
                aib19_ch0_x0y1, aib18_ch0_x0y1, aib17_ch0_x0y1,aib16_ch0_x0y1,
                aib15_ch0_x0y1, aib14_ch0_x0y1, aib13_ch0_x0y1,aib12_ch0_x0y1,
                aib11_ch0_x0y1, aib10_ch0_x0y1, aib9_ch0_x0y1, aib8_ch0_x0y1,
                aib7_ch0_x0y1,  aib6_ch0_x0y1,  aib5_ch0_x0y1, aib4_ch0_x0y1,
                aib3_ch0_x0y1,  aib2_ch0_x0y1,  aib1_ch0_x0y1, aib0_ch0_x0y1,
                aib19_ch0_x0y1, aib18_ch0_x0y1, aib17_ch0_x0y1,aib16_ch0_x0y1,
                aib15_ch0_x0y1, aib14_ch0_x0y1, aib13_ch0_x0y1,aib12_ch0_x0y1,
                aib11_ch0_x0y1, aib10_ch0_x0y1, aib9_ch0_x0y1, aib8_ch0_x0y1,
                aib7_ch0_x0y1,  aib6_ch0_x0y1,  aib5_ch0_x0y1, aib4_ch0_x0y1,
                aib3_ch0_x0y1,  aib2_ch0_x0y1,  aib1_ch0_x0y1, aib0_ch0_x0y1};

  assign AIB_CHAN7 = {aib95_ch1_x0y1, aib94_ch1_x0y1, 1'b1,          aib94_ch1_x0y1,
                aib91_ch1_x0y1, aib90_ch1_x0y1, aib89_ch1_x0y1,aib88_ch1_x0y1,
                aib87_ch1_x0y1, aib86_ch1_x0y1, aib85_ch1_x0y1,aib84_ch1_x0y1,
                aib85_ch1_x0y1, aib84_ch1_x0y1, aib81_ch1_x0y1,aib80_ch1_x0y1,
                aib79_ch1_x0y1, aib78_ch1_x0y1, aib77_ch1_x0y1,aib76_ch1_x0y1,
                aib75_ch1_x0y1, aib74_ch1_x0y1, aib73_ch1_x0y1,aib72_ch1_x0y1,
                aib71_ch1_x0y1, aib70_ch1_x0y1, aib69_ch1_x0y1,aib68_ch1_x0y1,
                aib67_ch1_x0y1, aib66_ch1_x0y1, 1'b1,          aib64_ch1_x0y1,
                aib63_ch1_x0y1, aib62_ch1_x0y1, 1'b1,          aib60_ch1_x0y1,
                aib59_ch1_x0y1, aib58_ch1_x0y1, aib57_ch1_x0y1,aib56_ch1_x0y1,
                aib55_ch1_x0y1, aib54_ch1_x0y1, aib53_ch1_x0y1,aib52_ch1_x0y1,
                aib51_ch1_x0y1, aib50_ch1_x0y1, aib49_ch1_x0y1,aib48_ch1_x0y1,
                aib47_ch1_x0y1, aib46_ch1_x0y1, aib45_ch1_x0y1,aib44_ch1_x0y1,
                aib41_ch1_x0y1, aib40_ch1_x0y1, aib41_ch1_x0y1,aib40_ch1_x0y1,
                aib19_ch1_x0y1, aib18_ch1_x0y1, aib17_ch1_x0y1,aib16_ch1_x0y1,
                aib15_ch1_x0y1, aib14_ch1_x0y1, aib13_ch1_x0y1,aib12_ch1_x0y1,
                aib11_ch1_x0y1, aib10_ch1_x0y1, aib9_ch1_x0y1, aib8_ch1_x0y1,
                aib7_ch1_x0y1,  aib6_ch1_x0y1,  aib5_ch1_x0y1, aib4_ch1_x0y1,
                aib3_ch1_x0y1,  aib2_ch1_x0y1,  aib1_ch1_x0y1, aib0_ch1_x0y1,
                aib19_ch1_x0y1, aib18_ch1_x0y1, aib17_ch1_x0y1,aib16_ch1_x0y1,
                aib15_ch1_x0y1, aib14_ch1_x0y1, aib13_ch1_x0y1,aib12_ch1_x0y1,
                aib11_ch1_x0y1, aib10_ch1_x0y1, aib9_ch1_x0y1, aib8_ch1_x0y1,
                aib7_ch1_x0y1,  aib6_ch1_x0y1,  aib5_ch1_x0y1, aib4_ch1_x0y1,
                aib3_ch1_x0y1,  aib2_ch1_x0y1,  aib1_ch1_x0y1, aib0_ch1_x0y1};

  assign AIB_CHAN8 = {aib95_ch2_x0y1, aib94_ch2_x0y1, 1'b1,          aib94_ch2_x0y1,
                aib91_ch2_x0y1, aib90_ch2_x0y1, aib89_ch2_x0y1,aib88_ch2_x0y1,
                aib87_ch2_x0y1, aib86_ch2_x0y1, aib85_ch2_x0y1,aib84_ch2_x0y1,
                aib85_ch2_x0y1, aib84_ch2_x0y1, aib81_ch2_x0y1,aib80_ch2_x0y1,
                aib79_ch2_x0y1, aib78_ch2_x0y1, aib77_ch2_x0y1,aib76_ch2_x0y1,
                aib75_ch2_x0y1, aib74_ch2_x0y1, aib73_ch2_x0y1,aib72_ch2_x0y1,
                aib71_ch2_x0y1, aib70_ch2_x0y1, aib69_ch2_x0y1,aib68_ch2_x0y1,
                aib67_ch2_x0y1, aib66_ch2_x0y1, 1'b1,          aib64_ch2_x0y1,
                aib63_ch2_x0y1, aib62_ch2_x0y1, 1'b1,          aib60_ch2_x0y1,
                aib59_ch2_x0y1, aib58_ch2_x0y1, aib57_ch2_x0y1,aib56_ch2_x0y1,
                aib55_ch2_x0y1, aib54_ch2_x0y1, aib53_ch2_x0y1,aib52_ch2_x0y1,
                aib51_ch2_x0y1, aib50_ch2_x0y1, aib49_ch2_x0y1,aib48_ch2_x0y1,
                aib47_ch2_x0y1, aib46_ch2_x0y1, aib45_ch2_x0y1,aib44_ch2_x0y1,
                aib41_ch2_x0y1, aib40_ch2_x0y1, aib41_ch2_x0y1,aib40_ch2_x0y1,
                aib19_ch2_x0y1, aib18_ch2_x0y1, aib17_ch2_x0y1,aib16_ch2_x0y1,
                aib15_ch2_x0y1, aib14_ch2_x0y1, aib13_ch2_x0y1,aib12_ch2_x0y1,
                aib11_ch2_x0y1, aib10_ch2_x0y1, aib9_ch2_x0y1, aib8_ch2_x0y1,
                aib7_ch2_x0y1,  aib6_ch2_x0y1,  aib5_ch2_x0y1, aib4_ch2_x0y1,
                aib3_ch2_x0y1,  aib2_ch2_x0y1,  aib1_ch2_x0y1, aib0_ch2_x0y1,
                aib19_ch2_x0y1, aib18_ch2_x0y1, aib17_ch2_x0y1,aib16_ch2_x0y1,
                aib15_ch2_x0y1, aib14_ch2_x0y1, aib13_ch2_x0y1,aib12_ch2_x0y1,
                aib11_ch2_x0y1, aib10_ch2_x0y1, aib9_ch2_x0y1, aib8_ch2_x0y1,
                aib7_ch2_x0y1,  aib6_ch2_x0y1,  aib5_ch2_x0y1, aib4_ch2_x0y1,
                aib3_ch2_x0y1,  aib2_ch2_x0y1,  aib1_ch2_x0y1, aib0_ch2_x0y1};

 assign AIB_CHAN9 = {aib95_ch3_x0y1, aib94_ch3_x0y1, 1'b1,          aib94_ch3_x0y1,
                aib91_ch3_x0y1, aib90_ch3_x0y1, aib89_ch3_x0y1,aib88_ch3_x0y1,
                aib87_ch3_x0y1, aib86_ch3_x0y1, aib85_ch3_x0y1,aib84_ch3_x0y1,
                aib85_ch3_x0y1, aib84_ch3_x0y1, aib81_ch3_x0y1,aib80_ch3_x0y1,
                aib79_ch3_x0y1, aib78_ch3_x0y1, aib77_ch3_x0y1,aib76_ch3_x0y1,
                aib75_ch3_x0y1, aib74_ch3_x0y1, aib73_ch3_x0y1,aib72_ch3_x0y1,
                aib71_ch3_x0y1, aib70_ch3_x0y1, aib69_ch3_x0y1,aib68_ch3_x0y1,
                aib67_ch3_x0y1, aib66_ch3_x0y1, 1'b1,          aib64_ch3_x0y1,
                aib63_ch3_x0y1, aib62_ch3_x0y1, 1'b1,          aib60_ch3_x0y1,
                aib59_ch3_x0y1, aib58_ch3_x0y1, aib57_ch3_x0y1,aib56_ch3_x0y1,
                aib55_ch3_x0y1, aib54_ch3_x0y1, aib53_ch3_x0y1,aib52_ch3_x0y1,
                aib51_ch3_x0y1, aib50_ch3_x0y1, aib49_ch3_x0y1,aib48_ch3_x0y1,
                aib47_ch3_x0y1, aib46_ch3_x0y1, aib45_ch3_x0y1,aib44_ch3_x0y1,
                aib41_ch3_x0y1, aib40_ch3_x0y1, aib41_ch3_x0y1,aib40_ch3_x0y1,
                aib19_ch3_x0y1, aib18_ch3_x0y1, aib17_ch3_x0y1,aib16_ch3_x0y1,
                aib15_ch3_x0y1, aib14_ch3_x0y1, aib13_ch3_x0y1,aib12_ch3_x0y1,
                aib11_ch3_x0y1, aib10_ch3_x0y1, aib9_ch3_x0y1, aib8_ch3_x0y1,
                aib7_ch3_x0y1,  aib6_ch3_x0y1,  aib5_ch3_x0y1, aib4_ch3_x0y1,
                aib3_ch3_x0y1,  aib2_ch3_x0y1,  aib1_ch3_x0y1, aib0_ch3_x0y1,
                aib19_ch3_x0y1, aib18_ch3_x0y1, aib17_ch3_x0y1,aib16_ch3_x0y1,
                aib15_ch3_x0y1, aib14_ch3_x0y1, aib13_ch3_x0y1,aib12_ch3_x0y1,
                aib11_ch3_x0y1, aib10_ch3_x0y1, aib9_ch3_x0y1, aib8_ch3_x0y1,
                aib7_ch3_x0y1,  aib6_ch3_x0y1,  aib5_ch3_x0y1, aib4_ch3_x0y1,
                aib3_ch3_x0y1,  aib2_ch3_x0y1,  aib1_ch3_x0y1, aib0_ch3_x0y1};

 assign AIB_CHAN10 = {aib95_ch4_x0y1, aib94_ch4_x0y1, 1'b1,         aib94_ch4_x0y1,
                aib91_ch4_x0y1, aib90_ch4_x0y1, aib89_ch4_x0y1,aib88_ch4_x0y1,
                aib87_ch4_x0y1, aib86_ch4_x0y1, aib85_ch4_x0y1,aib84_ch4_x0y1,
                aib85_ch4_x0y1, aib84_ch4_x0y1, aib81_ch4_x0y1,aib80_ch4_x0y1,
                aib79_ch4_x0y1, aib78_ch4_x0y1, aib77_ch4_x0y1,aib76_ch4_x0y1,
                aib75_ch4_x0y1, aib74_ch4_x0y1, aib73_ch4_x0y1,aib72_ch4_x0y1,
                aib71_ch4_x0y1, aib70_ch4_x0y1, aib69_ch4_x0y1,aib68_ch4_x0y1,
                aib67_ch4_x0y1, aib66_ch4_x0y1, 1'b1,          aib64_ch4_x0y1,
                aib63_ch4_x0y1, aib62_ch4_x0y1, 1'b1,          aib60_ch4_x0y1,
                aib59_ch4_x0y1, aib58_ch4_x0y1, aib57_ch4_x0y1,aib56_ch4_x0y1,
                aib55_ch4_x0y1, aib54_ch4_x0y1, aib53_ch4_x0y1,aib52_ch4_x0y1,
                aib51_ch4_x0y1, aib50_ch4_x0y1, aib49_ch4_x0y1,aib48_ch4_x0y1,
                aib47_ch4_x0y1, aib46_ch4_x0y1, aib45_ch4_x0y1,aib44_ch4_x0y1,
                aib41_ch4_x0y1, aib40_ch4_x0y1, aib41_ch4_x0y1,aib40_ch4_x0y1,
                aib19_ch4_x0y1, aib18_ch4_x0y1, aib17_ch4_x0y1,aib16_ch4_x0y1,
                aib15_ch4_x0y1, aib14_ch4_x0y1, aib13_ch4_x0y1,aib12_ch4_x0y1,
                aib11_ch4_x0y1, aib10_ch4_x0y1, aib9_ch4_x0y1, aib8_ch4_x0y1,
                aib7_ch4_x0y1,  aib6_ch4_x0y1,  aib5_ch4_x0y1, aib4_ch4_x0y1,
                aib3_ch4_x0y1,  aib2_ch4_x0y1,  aib1_ch4_x0y1, aib0_ch4_x0y1,
                aib19_ch4_x0y1, aib18_ch4_x0y1, aib17_ch4_x0y1,aib16_ch4_x0y1,
                aib15_ch4_x0y1, aib14_ch4_x0y1, aib13_ch4_x0y1,aib12_ch4_x0y1,
                aib11_ch4_x0y1, aib10_ch4_x0y1, aib9_ch4_x0y1, aib8_ch4_x0y1,
                aib7_ch4_x0y1,  aib6_ch4_x0y1,  aib5_ch4_x0y1, aib4_ch4_x0y1,
                aib3_ch4_x0y1,  aib2_ch4_x0y1,  aib1_ch4_x0y1, aib0_ch4_x0y1};

 assign AIB_CHAN11 = {aib95_ch5_x0y1, aib94_ch5_x0y1, 1'b1,         aib94_ch5_x0y1,
                aib91_ch5_x0y1, aib90_ch5_x0y1, aib89_ch5_x0y1,aib88_ch5_x0y1,
                aib87_ch5_x0y1, aib86_ch5_x0y1, aib85_ch5_x0y1,aib84_ch5_x0y1,
                aib85_ch5_x0y1, aib84_ch5_x0y1, aib81_ch5_x0y1,aib80_ch5_x0y1,
                aib79_ch5_x0y1, aib78_ch5_x0y1, aib77_ch5_x0y1,aib76_ch5_x0y1,
                aib75_ch5_x0y1, aib74_ch5_x0y1, aib73_ch5_x0y1,aib72_ch5_x0y1,
                aib71_ch5_x0y1, aib70_ch5_x0y1, aib69_ch5_x0y1,aib68_ch5_x0y1,
                aib67_ch5_x0y1, aib66_ch5_x0y1, 1'b1,          aib64_ch5_x0y1,
                aib63_ch5_x0y1, aib62_ch5_x0y1, 1'b1,          aib60_ch5_x0y1,
                aib59_ch5_x0y1, aib58_ch5_x0y1, aib57_ch5_x0y1,aib56_ch5_x0y1,
                aib55_ch5_x0y1, aib54_ch5_x0y1, aib53_ch5_x0y1,aib52_ch5_x0y1,
                aib51_ch5_x0y1, aib50_ch5_x0y1, aib49_ch5_x0y1,aib48_ch5_x0y1,
                aib47_ch5_x0y1, aib46_ch5_x0y1, aib45_ch5_x0y1,aib44_ch5_x0y1,
                aib41_ch5_x0y1, aib40_ch5_x0y1, aib41_ch5_x0y1,aib40_ch5_x0y1,
                aib19_ch5_x0y1, aib18_ch5_x0y1, aib17_ch5_x0y1,aib16_ch5_x0y1,
                aib15_ch5_x0y1, aib14_ch5_x0y1, aib13_ch5_x0y1,aib12_ch5_x0y1,
                aib11_ch5_x0y1, aib10_ch5_x0y1, aib9_ch5_x0y1, aib8_ch5_x0y1,
                aib7_ch5_x0y1,  aib6_ch5_x0y1,  aib5_ch5_x0y1, aib4_ch5_x0y1,
                aib3_ch5_x0y1,  aib2_ch5_x0y1,  aib1_ch5_x0y1, aib0_ch5_x0y1,
                aib19_ch5_x0y1, aib18_ch5_x0y1, aib17_ch5_x0y1,aib16_ch5_x0y1,
                aib15_ch5_x0y1, aib14_ch5_x0y1, aib13_ch5_x0y1,aib12_ch5_x0y1,
                aib11_ch5_x0y1, aib10_ch5_x0y1, aib9_ch5_x0y1, aib8_ch5_x0y1,
                aib7_ch5_x0y1,  aib6_ch5_x0y1,  aib5_ch5_x0y1, aib4_ch5_x0y1,
                aib3_ch5_x0y1,  aib2_ch5_x0y1,  aib1_ch5_x0y1, aib0_ch5_x0y1};

 assign AIB_CHAN12 = {aib95_ch0_x0y2, aib94_ch0_x0y2, 1'b1,         aib94_ch0_x0y2,
                aib91_ch0_x0y2, aib90_ch0_x0y2, aib89_ch0_x0y2,aib88_ch0_x0y2,
                aib87_ch0_x0y2, aib86_ch0_x0y2, aib85_ch0_x0y2,aib84_ch0_x0y2,
                aib85_ch0_x0y2, aib84_ch0_x0y2, aib81_ch0_x0y2,aib80_ch0_x0y2,
                aib79_ch0_x0y2, aib78_ch0_x0y2, aib77_ch0_x0y2,aib76_ch0_x0y2,
                aib75_ch0_x0y2, aib74_ch0_x0y2, aib73_ch0_x0y2,aib72_ch0_x0y2,
                aib71_ch0_x0y2, aib70_ch0_x0y2, aib69_ch0_x0y2,aib68_ch0_x0y2,
                aib67_ch0_x0y2, aib66_ch0_x0y2, 1'b1,          aib64_ch0_x0y2,
                aib63_ch0_x0y2, aib62_ch0_x0y2, 1'b1,          aib60_ch0_x0y2,
                aib59_ch0_x0y2, aib58_ch0_x0y2, aib57_ch0_x0y2,aib56_ch0_x0y2,
                aib55_ch0_x0y2, aib54_ch0_x0y2, aib53_ch0_x0y2,aib52_ch0_x0y2,
                aib51_ch0_x0y2, aib50_ch0_x0y2, aib49_ch0_x0y2,aib48_ch0_x0y2,
                aib47_ch0_x0y2, aib46_ch0_x0y2, aib45_ch0_x0y2,aib44_ch0_x0y2,
                aib41_ch0_x0y2, aib40_ch0_x0y2, aib41_ch0_x0y2,aib40_ch0_x0y2,
                aib19_ch0_x0y2, aib18_ch0_x0y2, aib17_ch0_x0y2,aib16_ch0_x0y2,
                aib15_ch0_x0y2, aib14_ch0_x0y2, aib13_ch0_x0y2,aib12_ch0_x0y2,
                aib11_ch0_x0y2, aib10_ch0_x0y2, aib9_ch0_x0y2, aib8_ch0_x0y2,
                aib7_ch0_x0y2,  aib6_ch0_x0y2,  aib5_ch0_x0y2, aib4_ch0_x0y2,
                aib3_ch0_x0y2,  aib2_ch0_x0y2,  aib1_ch0_x0y2, aib0_ch0_x0y2,
                aib19_ch0_x0y2, aib18_ch0_x0y2, aib17_ch0_x0y2,aib16_ch0_x0y2,
                aib15_ch0_x0y2, aib14_ch0_x0y2, aib13_ch0_x0y2,aib12_ch0_x0y2,
                aib11_ch0_x0y2, aib10_ch0_x0y2, aib9_ch0_x0y2, aib8_ch0_x0y2,
                aib7_ch0_x0y2,  aib6_ch0_x0y2,  aib5_ch0_x0y2, aib4_ch0_x0y2,
                aib3_ch0_x0y2,  aib2_ch0_x0y2,  aib1_ch0_x0y2, aib0_ch0_x0y2};

 assign  AIB_CHAN13 = {aib95_ch1_x0y2, aib94_ch1_x0y2, 1'b1,         aib94_ch1_x0y2,
                aib91_ch1_x0y2, aib90_ch1_x0y2, aib89_ch1_x0y2,aib88_ch1_x0y2,
                aib87_ch1_x0y2, aib86_ch1_x0y2, aib85_ch1_x0y2,aib84_ch1_x0y2,
                aib85_ch1_x0y2, aib84_ch1_x0y2, aib81_ch1_x0y2,aib80_ch1_x0y2,
                aib79_ch1_x0y2, aib78_ch1_x0y2, aib77_ch1_x0y2,aib76_ch1_x0y2,
                aib75_ch1_x0y2, aib74_ch1_x0y2, aib73_ch1_x0y2,aib72_ch1_x0y2,
                aib71_ch1_x0y2, aib70_ch1_x0y2, aib69_ch1_x0y2,aib68_ch1_x0y2,
                aib67_ch1_x0y2, aib66_ch1_x0y2, 1'b1,          aib64_ch1_x0y2,
                aib63_ch1_x0y2, aib62_ch1_x0y2, 1'b1,          aib60_ch1_x0y2,
                aib59_ch1_x0y2, aib58_ch1_x0y2, aib57_ch1_x0y2,aib56_ch1_x0y2,
                aib55_ch1_x0y2, aib54_ch1_x0y2, aib53_ch1_x0y2,aib52_ch1_x0y2,
                aib51_ch1_x0y2, aib50_ch1_x0y2, aib49_ch1_x0y2,aib48_ch1_x0y2,
                aib47_ch1_x0y2, aib46_ch1_x0y2, aib45_ch1_x0y2,aib44_ch1_x0y2,
                aib41_ch1_x0y2, aib40_ch1_x0y2, aib41_ch1_x0y2,aib40_ch1_x0y2,
                aib19_ch1_x0y2, aib18_ch1_x0y2, aib17_ch1_x0y2,aib16_ch1_x0y2,
                aib15_ch1_x0y2, aib14_ch1_x0y2, aib13_ch1_x0y2,aib12_ch1_x0y2,
                aib11_ch1_x0y2, aib10_ch1_x0y2, aib9_ch1_x0y2, aib8_ch1_x0y2,
                aib7_ch1_x0y2,  aib6_ch1_x0y2,  aib5_ch1_x0y2, aib4_ch1_x0y2,
                aib3_ch1_x0y2,  aib2_ch1_x0y2,  aib1_ch1_x0y2, aib0_ch1_x0y2,
                aib19_ch1_x0y2, aib18_ch1_x0y2, aib17_ch1_x0y2,aib16_ch1_x0y2,
                aib15_ch1_x0y2, aib14_ch1_x0y2, aib13_ch1_x0y2,aib12_ch1_x0y2,
                aib11_ch1_x0y2, aib10_ch1_x0y2, aib9_ch1_x0y2, aib8_ch1_x0y2,
                aib7_ch1_x0y2,  aib6_ch1_x0y2,  aib5_ch1_x0y2, aib4_ch1_x0y2,
                aib3_ch1_x0y2,  aib2_ch1_x0y2,  aib1_ch1_x0y2, aib0_ch1_x0y2};

 assign AIB_CHAN14 ={aib95_ch2_x0y2, aib94_ch2_x0y2, 1'b1,         aib94_ch2_x0y2,
                aib91_ch2_x0y2, aib90_ch2_x0y2, aib89_ch2_x0y2,aib88_ch2_x0y2,
                aib87_ch2_x0y2, aib86_ch2_x0y2, aib85_ch2_x0y2,aib84_ch2_x0y2,
                aib85_ch2_x0y2, aib84_ch2_x0y2, aib81_ch2_x0y2,aib80_ch2_x0y2,
                aib79_ch2_x0y2, aib78_ch2_x0y2, aib77_ch2_x0y2,aib76_ch2_x0y2,
                aib75_ch2_x0y2, aib74_ch2_x0y2, aib73_ch2_x0y2,aib72_ch2_x0y2,
                aib71_ch2_x0y2, aib70_ch2_x0y2, aib69_ch2_x0y2,aib68_ch2_x0y2,
                aib67_ch2_x0y2, aib66_ch2_x0y2, 1'b1,          aib64_ch2_x0y2,
                aib63_ch2_x0y2, aib62_ch2_x0y2, 1'b1,          aib60_ch2_x0y2,
                aib59_ch2_x0y2, aib58_ch2_x0y2, aib57_ch2_x0y2,aib56_ch2_x0y2,
                aib55_ch2_x0y2, aib54_ch2_x0y2, aib53_ch2_x0y2,aib52_ch2_x0y2,
                aib51_ch2_x0y2, aib50_ch2_x0y2, aib49_ch2_x0y2,aib48_ch2_x0y2,
                aib47_ch2_x0y2, aib46_ch2_x0y2, aib45_ch2_x0y2,aib44_ch2_x0y2,
                aib41_ch2_x0y2, aib40_ch2_x0y2, aib41_ch2_x0y2,aib40_ch2_x0y2,
                aib19_ch2_x0y2, aib18_ch2_x0y2, aib17_ch2_x0y2,aib16_ch2_x0y2,
                aib15_ch2_x0y2, aib14_ch2_x0y2, aib13_ch2_x0y2,aib12_ch2_x0y2,
                aib11_ch2_x0y2, aib10_ch2_x0y2, aib9_ch2_x0y2, aib8_ch2_x0y2,
                aib7_ch2_x0y2,  aib6_ch2_x0y2,  aib5_ch2_x0y2, aib4_ch2_x0y2,
                aib3_ch2_x0y2,  aib2_ch2_x0y2,  aib1_ch2_x0y2, aib0_ch2_x0y2,
                aib19_ch2_x0y2, aib18_ch2_x0y2, aib17_ch2_x0y2,aib16_ch2_x0y2,
                aib15_ch2_x0y2, aib14_ch2_x0y2, aib13_ch2_x0y2,aib12_ch2_x0y2,
                aib11_ch2_x0y2, aib10_ch2_x0y2, aib9_ch2_x0y2, aib8_ch2_x0y2,
                aib7_ch2_x0y2,  aib6_ch2_x0y2,  aib5_ch2_x0y2, aib4_ch2_x0y2,
                aib3_ch2_x0y2,  aib2_ch2_x0y2,  aib1_ch2_x0y2, aib0_ch2_x0y2};

  assign  AIB_CHAN15 = {aib95_ch3_x0y2, aib94_ch3_x0y2, 1'b1,         aib94_ch3_x0y2,
                aib91_ch3_x0y2, aib90_ch3_x0y2, aib89_ch3_x0y2,aib88_ch3_x0y2,
                aib87_ch3_x0y2, aib86_ch3_x0y2, aib85_ch3_x0y2,aib84_ch3_x0y2,
                aib85_ch3_x0y2, aib84_ch3_x0y2, aib81_ch3_x0y2,aib80_ch3_x0y2,
                aib79_ch3_x0y2, aib78_ch3_x0y2, aib77_ch3_x0y2,aib76_ch3_x0y2,
                aib75_ch3_x0y2, aib74_ch3_x0y2, aib73_ch3_x0y2,aib72_ch3_x0y2,
                aib71_ch3_x0y2, aib70_ch3_x0y2, aib69_ch3_x0y2,aib68_ch3_x0y2,
                aib67_ch3_x0y2, aib66_ch3_x0y2, 1'b1,          aib64_ch3_x0y2,
                aib63_ch3_x0y2, aib62_ch3_x0y2, 1'b1,          aib60_ch3_x0y2,
                aib59_ch3_x0y2, aib58_ch3_x0y2, aib57_ch3_x0y2,aib56_ch3_x0y2,
                aib55_ch3_x0y2, aib54_ch3_x0y2, aib53_ch3_x0y2,aib52_ch3_x0y2,
                aib51_ch3_x0y2, aib50_ch3_x0y2, aib49_ch3_x0y2,aib48_ch3_x0y2,
                aib47_ch3_x0y2, aib46_ch3_x0y2, aib45_ch3_x0y2,aib44_ch3_x0y2,
                aib41_ch3_x0y2, aib40_ch3_x0y2, aib41_ch3_x0y2,aib40_ch3_x0y2,
                aib19_ch3_x0y2, aib18_ch3_x0y2, aib17_ch3_x0y2,aib16_ch3_x0y2,
                aib15_ch3_x0y2, aib14_ch3_x0y2, aib13_ch3_x0y2,aib12_ch3_x0y2,
                aib11_ch3_x0y2, aib10_ch3_x0y2, aib9_ch3_x0y2, aib8_ch3_x0y2,
                aib7_ch3_x0y2,  aib6_ch3_x0y2,  aib5_ch3_x0y2, aib4_ch3_x0y2,
                aib3_ch3_x0y2,  aib2_ch3_x0y2,  aib1_ch3_x0y2, aib0_ch3_x0y2,
                aib19_ch3_x0y2, aib18_ch3_x0y2, aib17_ch3_x0y2,aib16_ch3_x0y2,
                aib15_ch3_x0y2, aib14_ch3_x0y2, aib13_ch3_x0y2,aib12_ch3_x0y2,
                aib11_ch3_x0y2, aib10_ch3_x0y2, aib9_ch3_x0y2, aib8_ch3_x0y2,
                aib7_ch3_x0y2,  aib6_ch3_x0y2,  aib5_ch3_x0y2, aib4_ch3_x0y2,
                aib3_ch3_x0y2,  aib2_ch3_x0y2,  aib1_ch3_x0y2, aib0_ch3_x0y2};

 assign AIB_CHAN16 = {aib95_ch4_x0y2, aib94_ch4_x0y2, 1'b1,         aib94_ch4_x0y2,
                aib91_ch4_x0y2, aib90_ch4_x0y2, aib89_ch4_x0y2,aib88_ch4_x0y2,
                aib87_ch4_x0y2, aib86_ch4_x0y2, aib85_ch4_x0y2,aib84_ch4_x0y2,
                aib85_ch4_x0y2, aib84_ch4_x0y2, aib81_ch4_x0y2,aib80_ch4_x0y2,
                aib79_ch4_x0y2, aib78_ch4_x0y2, aib77_ch4_x0y2,aib76_ch4_x0y2,
                aib75_ch4_x0y2, aib74_ch4_x0y2, aib73_ch4_x0y2,aib72_ch4_x0y2,
                aib71_ch4_x0y2, aib70_ch4_x0y2, aib69_ch4_x0y2,aib68_ch4_x0y2,
                aib67_ch4_x0y2, aib66_ch4_x0y2, 1'b1,          aib64_ch4_x0y2,
                aib63_ch4_x0y2, aib62_ch4_x0y2, 1'b1,          aib60_ch4_x0y2,
                aib59_ch4_x0y2, aib58_ch4_x0y2, aib57_ch4_x0y2,aib56_ch4_x0y2,
                aib55_ch4_x0y2, aib54_ch4_x0y2, aib53_ch4_x0y2,aib52_ch4_x0y2,
                aib51_ch4_x0y2, aib50_ch4_x0y2, aib49_ch4_x0y2,aib48_ch4_x0y2,
                aib47_ch4_x0y2, aib46_ch4_x0y2, aib45_ch4_x0y2,aib44_ch4_x0y2,
                aib41_ch4_x0y2, aib40_ch4_x0y2, aib41_ch4_x0y2,aib40_ch4_x0y2,
                aib19_ch4_x0y2, aib18_ch4_x0y2, aib17_ch4_x0y2,aib16_ch4_x0y2,
                aib15_ch4_x0y2, aib14_ch4_x0y2, aib13_ch4_x0y2,aib12_ch4_x0y2,
                aib11_ch4_x0y2, aib10_ch4_x0y2, aib9_ch4_x0y2, aib8_ch4_x0y2,
                aib7_ch4_x0y2,  aib6_ch4_x0y2,  aib5_ch4_x0y2, aib4_ch4_x0y2,
                aib3_ch4_x0y2,  aib2_ch4_x0y2,  aib1_ch4_x0y2, aib0_ch4_x0y2,
                aib19_ch4_x0y2, aib18_ch4_x0y2, aib17_ch4_x0y2,aib16_ch4_x0y2,
                aib15_ch4_x0y2, aib14_ch4_x0y2, aib13_ch4_x0y2,aib12_ch4_x0y2,
                aib11_ch4_x0y2, aib10_ch4_x0y2, aib9_ch4_x0y2, aib8_ch4_x0y2,
                aib7_ch4_x0y2,  aib6_ch4_x0y2,  aib5_ch4_x0y2, aib4_ch4_x0y2,
                aib3_ch4_x0y2,  aib2_ch4_x0y2,  aib1_ch4_x0y2, aib0_ch4_x0y2};

  assign AIB_CHAN17 = {aib95_ch5_x0y2, aib94_ch5_x0y2, 1'b1,         aib94_ch5_x0y2,
                aib91_ch5_x0y2, aib90_ch5_x0y2, aib89_ch5_x0y2,aib88_ch5_x0y2,
                aib87_ch5_x0y2, aib86_ch5_x0y2, aib85_ch5_x0y2,aib84_ch5_x0y2,
                aib85_ch5_x0y2, aib84_ch5_x0y2, aib81_ch5_x0y2,aib80_ch5_x0y2,
                aib79_ch5_x0y2, aib78_ch5_x0y2, aib77_ch5_x0y2,aib76_ch5_x0y2,
                aib75_ch5_x0y2, aib74_ch5_x0y2, aib73_ch5_x0y2,aib72_ch5_x0y2,
                aib71_ch5_x0y2, aib70_ch5_x0y2, aib69_ch5_x0y2,aib68_ch5_x0y2,
                aib67_ch5_x0y2, aib66_ch5_x0y2, 1'b1,          aib64_ch5_x0y2,
                aib63_ch5_x0y2, aib62_ch5_x0y2, 1'b1,          aib60_ch5_x0y2,
                aib59_ch5_x0y2, aib58_ch5_x0y2, aib57_ch5_x0y2,aib56_ch5_x0y2,
                aib55_ch5_x0y2, aib54_ch5_x0y2, aib53_ch5_x0y2,aib52_ch5_x0y2,
                aib51_ch5_x0y2, aib50_ch5_x0y2, aib49_ch5_x0y2,aib48_ch5_x0y2,
                aib47_ch5_x0y2, aib46_ch5_x0y2, aib45_ch5_x0y2,aib44_ch5_x0y2,
                aib41_ch5_x0y2, aib40_ch5_x0y2, aib41_ch5_x0y2,aib40_ch5_x0y2,
                aib19_ch5_x0y2, aib18_ch5_x0y2, aib17_ch5_x0y2,aib16_ch5_x0y2,
                aib15_ch5_x0y2, aib14_ch5_x0y2, aib13_ch5_x0y2,aib12_ch5_x0y2,
                aib11_ch5_x0y2, aib10_ch5_x0y2, aib9_ch5_x0y2, aib8_ch5_x0y2,
                aib7_ch5_x0y2,  aib6_ch5_x0y2,  aib5_ch5_x0y2, aib4_ch5_x0y2,
                aib3_ch5_x0y2,  aib2_ch5_x0y2,  aib1_ch5_x0y2, aib0_ch5_x0y2,
                aib19_ch5_x0y2, aib18_ch5_x0y2, aib17_ch5_x0y2,aib16_ch5_x0y2,
                aib15_ch5_x0y2, aib14_ch5_x0y2, aib13_ch5_x0y2,aib12_ch5_x0y2,
                aib11_ch5_x0y2, aib10_ch5_x0y2, aib9_ch5_x0y2, aib8_ch5_x0y2,
                aib7_ch5_x0y2,  aib6_ch5_x0y2,  aib5_ch5_x0y2, aib4_ch5_x0y2,
                aib3_ch5_x0y2,  aib2_ch5_x0y2,  aib1_ch5_x0y2, aib0_ch5_x0y2};

 assign AIB_CHAN18 = {aib95_ch0_x0y3, aib94_ch0_x0y3, 1'b1,         aib94_ch0_x0y3,
                aib91_ch0_x0y3, aib90_ch0_x0y3, aib89_ch0_x0y3,aib88_ch0_x0y3,
                aib87_ch0_x0y3, aib86_ch0_x0y3, aib85_ch0_x0y3,aib84_ch0_x0y3,
                aib85_ch0_x0y3, aib84_ch0_x0y3, aib81_ch0_x0y3,aib80_ch0_x0y3,
                aib79_ch0_x0y3, aib78_ch0_x0y3, aib77_ch0_x0y3,aib76_ch0_x0y3,
                aib75_ch0_x0y3, aib74_ch0_x0y3, aib73_ch0_x0y3,aib72_ch0_x0y3,
                aib71_ch0_x0y3, aib70_ch0_x0y3, aib69_ch0_x0y3,aib68_ch0_x0y3,
                aib67_ch0_x0y3, aib66_ch0_x0y3, 1'b1,          aib64_ch0_x0y3,
                aib63_ch0_x0y3, aib62_ch0_x0y3, 1'b1,          aib60_ch0_x0y3,
                aib59_ch0_x0y3, aib58_ch0_x0y3, aib57_ch0_x0y3,aib56_ch0_x0y3,
                aib55_ch0_x0y3, aib54_ch0_x0y3, aib53_ch0_x0y3,aib52_ch0_x0y3,
                aib51_ch0_x0y3, aib50_ch0_x0y3, aib49_ch0_x0y3,aib48_ch0_x0y3,
                aib47_ch0_x0y3, aib46_ch0_x0y3, aib45_ch0_x0y3,aib44_ch0_x0y3,
                aib41_ch0_x0y3, aib40_ch0_x0y3, aib41_ch0_x0y3,aib40_ch0_x0y3,
                aib19_ch0_x0y3, aib18_ch0_x0y3, aib17_ch0_x0y3,aib16_ch0_x0y3,
                aib15_ch0_x0y3, aib14_ch0_x0y3, aib13_ch0_x0y3,aib12_ch0_x0y3,
                aib11_ch0_x0y3, aib10_ch0_x0y3, aib9_ch0_x0y3, aib8_ch0_x0y3,
                aib7_ch0_x0y3,  aib6_ch0_x0y3,  aib5_ch0_x0y3, aib4_ch0_x0y3,
                aib3_ch0_x0y3,  aib2_ch0_x0y3,  aib1_ch0_x0y3, aib0_ch0_x0y3,
                aib19_ch0_x0y3, aib18_ch0_x0y3, aib17_ch0_x0y3,aib16_ch0_x0y3,
                aib15_ch0_x0y3, aib14_ch0_x0y3, aib13_ch0_x0y3,aib12_ch0_x0y3,
                aib11_ch0_x0y3, aib10_ch0_x0y3, aib9_ch0_x0y3, aib8_ch0_x0y3,
                aib7_ch0_x0y3,  aib6_ch0_x0y3,  aib5_ch0_x0y3, aib4_ch0_x0y3,
                aib3_ch0_x0y3,  aib2_ch0_x0y3,  aib1_ch0_x0y3, aib0_ch0_x0y3};

 assign AIB_CHAN19 = {aib95_ch1_x0y3, aib94_ch1_x0y3, 1'b1,         aib94_ch1_x0y3,
                aib91_ch1_x0y3, aib90_ch1_x0y3, aib89_ch1_x0y3,aib88_ch1_x0y3,
                aib87_ch1_x0y3, aib86_ch1_x0y3, aib85_ch1_x0y3,aib84_ch1_x0y3,
                aib85_ch1_x0y3, aib84_ch1_x0y3, aib81_ch1_x0y3,aib80_ch1_x0y3,
                aib79_ch1_x0y3, aib78_ch1_x0y3, aib77_ch1_x0y3,aib76_ch1_x0y3,
                aib75_ch1_x0y3, aib74_ch1_x0y3, aib73_ch1_x0y3,aib72_ch1_x0y3,
                aib71_ch1_x0y3, aib70_ch1_x0y3, aib69_ch1_x0y3,aib68_ch1_x0y3,
                aib67_ch1_x0y3, aib66_ch1_x0y3, 1'b1,          aib64_ch1_x0y3,
                aib63_ch1_x0y3, aib62_ch1_x0y3, 1'b1,          aib60_ch1_x0y3,
                aib59_ch1_x0y3, aib58_ch1_x0y3, aib57_ch1_x0y3,aib56_ch1_x0y3,
                aib55_ch1_x0y3, aib54_ch1_x0y3, aib53_ch1_x0y3,aib52_ch1_x0y3,
                aib51_ch1_x0y3, aib50_ch1_x0y3, aib49_ch1_x0y3,aib48_ch1_x0y3,
                aib47_ch1_x0y3, aib46_ch1_x0y3, aib45_ch1_x0y3,aib44_ch1_x0y3,
                aib41_ch1_x0y3, aib40_ch1_x0y3, aib41_ch1_x0y3,aib40_ch1_x0y3,
                aib19_ch1_x0y3, aib18_ch1_x0y3, aib17_ch1_x0y3,aib16_ch1_x0y3,
                aib15_ch1_x0y3, aib14_ch1_x0y3, aib13_ch1_x0y3,aib12_ch1_x0y3,
                aib11_ch1_x0y3, aib10_ch1_x0y3, aib9_ch1_x0y3, aib8_ch1_x0y3,
                aib7_ch1_x0y3,  aib6_ch1_x0y3,  aib5_ch1_x0y3, aib4_ch1_x0y3,
                aib3_ch1_x0y3,  aib2_ch1_x0y3,  aib1_ch1_x0y3, aib0_ch1_x0y3,
                aib19_ch1_x0y3, aib18_ch1_x0y3, aib17_ch1_x0y3,aib16_ch1_x0y3,
                aib15_ch1_x0y3, aib14_ch1_x0y3, aib13_ch1_x0y3,aib12_ch1_x0y3,
                aib11_ch1_x0y3, aib10_ch1_x0y3, aib9_ch1_x0y3, aib8_ch1_x0y3,
                aib7_ch1_x0y3,  aib6_ch1_x0y3,  aib5_ch1_x0y3, aib4_ch1_x0y3,
                aib3_ch1_x0y3,  aib2_ch1_x0y3,  aib1_ch1_x0y3, aib0_ch1_x0y3};

 assign AIB_CHAN20 = {aib95_ch2_x0y3, aib94_ch2_x0y3, 1'b1,         aib94_ch2_x0y3,
                aib91_ch2_x0y3, aib90_ch2_x0y3, aib89_ch2_x0y3,aib88_ch2_x0y3,
                aib87_ch2_x0y3, aib86_ch2_x0y3, aib85_ch2_x0y3,aib84_ch2_x0y3,
                aib85_ch2_x0y3, aib84_ch2_x0y3, aib81_ch2_x0y3,aib80_ch2_x0y3,
                aib79_ch2_x0y3, aib78_ch2_x0y3, aib77_ch2_x0y3,aib76_ch2_x0y3,
                aib75_ch2_x0y3, aib74_ch2_x0y3, aib73_ch2_x0y3,aib72_ch2_x0y3,
                aib71_ch2_x0y3, aib70_ch2_x0y3, aib69_ch2_x0y3,aib68_ch2_x0y3,
                aib67_ch2_x0y3, aib66_ch2_x0y3, 1'b1,          aib64_ch2_x0y3,
                aib63_ch2_x0y3, aib62_ch2_x0y3, 1'b1,          aib60_ch2_x0y3,
                aib59_ch2_x0y3, aib58_ch2_x0y3, aib57_ch2_x0y3,aib56_ch2_x0y3,
                aib55_ch2_x0y3, aib54_ch2_x0y3, aib53_ch2_x0y3,aib52_ch2_x0y3,
                aib51_ch2_x0y3, aib50_ch2_x0y3, aib49_ch2_x0y3,aib48_ch2_x0y3,
                aib47_ch2_x0y3, aib46_ch2_x0y3, aib45_ch2_x0y3,aib44_ch2_x0y3,
                aib41_ch2_x0y3, aib40_ch2_x0y3, aib41_ch2_x0y3,aib40_ch2_x0y3,
                aib19_ch2_x0y3, aib18_ch2_x0y3, aib17_ch2_x0y3,aib16_ch2_x0y3,
                aib15_ch2_x0y3, aib14_ch2_x0y3, aib13_ch2_x0y3,aib12_ch2_x0y3,
                aib11_ch2_x0y3, aib10_ch2_x0y3, aib9_ch2_x0y3, aib8_ch2_x0y3,
                aib7_ch2_x0y3,  aib6_ch2_x0y3,  aib5_ch2_x0y3, aib4_ch2_x0y3,
                aib3_ch2_x0y3,  aib2_ch2_x0y3,  aib1_ch2_x0y3, aib0_ch2_x0y3,
                aib19_ch2_x0y3, aib18_ch2_x0y3, aib17_ch2_x0y3,aib16_ch2_x0y3,
                aib15_ch2_x0y3, aib14_ch2_x0y3, aib13_ch2_x0y3,aib12_ch2_x0y3,
                aib11_ch2_x0y3, aib10_ch2_x0y3, aib9_ch2_x0y3, aib8_ch2_x0y3,
                aib7_ch2_x0y3,  aib6_ch2_x0y3,  aib5_ch2_x0y3, aib4_ch2_x0y3,
                aib3_ch2_x0y3,  aib2_ch2_x0y3,  aib1_ch2_x0y3, aib0_ch2_x0y3};

 assign AIB_CHAN21 = {aib95_ch3_x0y3, aib94_ch3_x0y3, 1'b1,         aib94_ch3_x0y3,
                aib91_ch3_x0y3, aib90_ch3_x0y3, aib89_ch3_x0y3,aib88_ch3_x0y3,
                aib87_ch3_x0y3, aib86_ch3_x0y3, aib85_ch3_x0y3,aib84_ch3_x0y3,
                aib85_ch3_x0y3, aib84_ch3_x0y3, aib81_ch3_x0y3,aib80_ch3_x0y3,
                aib79_ch3_x0y3, aib78_ch3_x0y3, aib77_ch3_x0y3,aib76_ch3_x0y3,
                aib75_ch3_x0y3, aib74_ch3_x0y3, aib73_ch3_x0y3,aib72_ch3_x0y3,
                aib71_ch3_x0y3, aib70_ch3_x0y3, aib69_ch3_x0y3,aib68_ch3_x0y3,
                aib67_ch3_x0y3, aib66_ch3_x0y3, 1'b1,          aib64_ch3_x0y3,
                aib63_ch3_x0y3, aib62_ch3_x0y3, 1'b1,          aib60_ch3_x0y3,
                aib59_ch3_x0y3, aib58_ch3_x0y3, aib57_ch3_x0y3,aib56_ch3_x0y3,
                aib55_ch3_x0y3, aib54_ch3_x0y3, aib53_ch3_x0y3,aib52_ch3_x0y3,
                aib51_ch3_x0y3, aib50_ch3_x0y3, aib49_ch3_x0y3,aib48_ch3_x0y3,
                aib47_ch3_x0y3, aib46_ch3_x0y3, aib45_ch3_x0y3,aib44_ch3_x0y3,
                aib41_ch3_x0y3, aib40_ch3_x0y3, aib41_ch3_x0y3,aib40_ch3_x0y3,
                aib19_ch3_x0y3, aib18_ch3_x0y3, aib17_ch3_x0y3,aib16_ch3_x0y3,
                aib15_ch3_x0y3, aib14_ch3_x0y3, aib13_ch3_x0y3,aib12_ch3_x0y3,
                aib11_ch3_x0y3, aib10_ch3_x0y3, aib9_ch3_x0y3, aib8_ch3_x0y3,
                aib7_ch3_x0y3,  aib6_ch3_x0y3,  aib5_ch3_x0y3, aib4_ch3_x0y3,
                aib3_ch3_x0y3,  aib2_ch3_x0y3,  aib1_ch3_x0y3, aib0_ch3_x0y3,
                aib19_ch3_x0y3, aib18_ch3_x0y3, aib17_ch3_x0y3,aib16_ch3_x0y3,
                aib15_ch3_x0y3, aib14_ch3_x0y3, aib13_ch3_x0y3,aib12_ch3_x0y3,
                aib11_ch3_x0y3, aib10_ch3_x0y3, aib9_ch3_x0y3, aib8_ch3_x0y3,
                aib7_ch3_x0y3,  aib6_ch3_x0y3,  aib5_ch3_x0y3, aib4_ch3_x0y3,
                aib3_ch3_x0y3,  aib2_ch3_x0y3,  aib1_ch3_x0y3, aib0_ch3_x0y3};

 assign AIB_CHAN22 = {aib95_ch4_x0y3, aib94_ch4_x0y3, 1'b1,         aib94_ch4_x0y3,
                aib91_ch4_x0y3, aib90_ch4_x0y3, aib89_ch4_x0y3,aib88_ch4_x0y3,
                aib87_ch4_x0y3, aib86_ch4_x0y3, aib85_ch4_x0y3,aib84_ch4_x0y3,
                aib85_ch4_x0y3, aib84_ch4_x0y3, aib81_ch4_x0y3,aib80_ch4_x0y3,
                aib79_ch4_x0y3, aib78_ch4_x0y3, aib77_ch4_x0y3,aib76_ch4_x0y3,
                aib75_ch4_x0y3, aib74_ch4_x0y3, aib73_ch4_x0y3,aib72_ch4_x0y3,
                aib71_ch4_x0y3, aib70_ch4_x0y3, aib69_ch4_x0y3,aib68_ch4_x0y3,
                aib67_ch4_x0y3, aib66_ch4_x0y3, 1'b1,          aib64_ch4_x0y3,
                aib63_ch4_x0y3, aib62_ch4_x0y3, 1'b1,          aib60_ch4_x0y3,
                aib59_ch4_x0y3, aib58_ch4_x0y3, aib57_ch4_x0y3,aib56_ch4_x0y3,
                aib55_ch4_x0y3, aib54_ch4_x0y3, aib53_ch4_x0y3,aib52_ch4_x0y3,
                aib51_ch4_x0y3, aib50_ch4_x0y3, aib49_ch4_x0y3,aib48_ch4_x0y3,
                aib47_ch4_x0y3, aib46_ch4_x0y3, aib45_ch4_x0y3,aib44_ch4_x0y3,
                aib41_ch4_x0y3, aib40_ch4_x0y3, aib41_ch4_x0y3,aib40_ch4_x0y3,
                aib19_ch4_x0y3, aib18_ch4_x0y3, aib17_ch4_x0y3,aib16_ch4_x0y3,
                aib15_ch4_x0y3, aib14_ch4_x0y3, aib13_ch4_x0y3,aib12_ch4_x0y3,
                aib11_ch4_x0y3, aib10_ch4_x0y3, aib9_ch4_x0y3, aib8_ch4_x0y3,
                aib7_ch4_x0y3,  aib6_ch4_x0y3,  aib5_ch4_x0y3, aib4_ch4_x0y3,
                aib3_ch4_x0y3,  aib2_ch4_x0y3,  aib1_ch4_x0y3, aib0_ch4_x0y3,
                aib19_ch4_x0y3, aib18_ch4_x0y3, aib17_ch4_x0y3,aib16_ch4_x0y3,
                aib15_ch4_x0y3, aib14_ch4_x0y3, aib13_ch4_x0y3,aib12_ch4_x0y3,
                aib11_ch4_x0y3, aib10_ch4_x0y3, aib9_ch4_x0y3, aib8_ch4_x0y3,
                aib7_ch4_x0y3,  aib6_ch4_x0y3,  aib5_ch4_x0y3, aib4_ch4_x0y3,
                aib3_ch4_x0y3,  aib2_ch4_x0y3,  aib1_ch4_x0y3, aib0_ch4_x0y3};

 assign AIB_CHAN23 = {aib95_ch5_x0y3, aib94_ch5_x0y3, 1'b1,         aib94_ch5_x0y3,
                aib91_ch5_x0y3, aib90_ch5_x0y3, aib89_ch5_x0y3,aib88_ch5_x0y3,
                aib87_ch5_x0y3, aib86_ch5_x0y3, aib85_ch5_x0y3,aib84_ch5_x0y3,
                aib85_ch5_x0y3, aib84_ch5_x0y3, aib81_ch5_x0y3,aib80_ch5_x0y3,
                aib79_ch5_x0y3, aib78_ch5_x0y3, aib77_ch5_x0y3,aib76_ch5_x0y3,
                aib75_ch5_x0y3, aib74_ch5_x0y3, aib73_ch5_x0y3,aib72_ch5_x0y3,
                aib71_ch5_x0y3, aib70_ch5_x0y3, aib69_ch5_x0y3,aib68_ch5_x0y3,
                aib67_ch5_x0y3, aib66_ch5_x0y3, 1'b1,          aib64_ch5_x0y3,
                aib63_ch5_x0y3, aib62_ch5_x0y3, 1'b1,          aib60_ch5_x0y3,
                aib59_ch5_x0y3, aib58_ch5_x0y3, aib57_ch5_x0y3,aib56_ch5_x0y3,
                aib55_ch5_x0y3, aib54_ch5_x0y3, aib53_ch5_x0y3,aib52_ch5_x0y3,
                aib51_ch5_x0y3, aib50_ch5_x0y3, aib49_ch5_x0y3,aib48_ch5_x0y3,
                aib47_ch5_x0y3, aib46_ch5_x0y3, aib45_ch5_x0y3,aib44_ch5_x0y3,
                aib41_ch5_x0y3, aib40_ch5_x0y3, aib41_ch5_x0y3,aib40_ch5_x0y3,
                aib19_ch5_x0y3, aib18_ch5_x0y3, aib17_ch5_x0y3,aib16_ch5_x0y3,
                aib15_ch5_x0y3, aib14_ch5_x0y3, aib13_ch5_x0y3,aib12_ch5_x0y3,
                aib11_ch5_x0y3, aib10_ch5_x0y3, aib9_ch5_x0y3, aib8_ch5_x0y3,
                aib7_ch5_x0y3,  aib6_ch5_x0y3,  aib5_ch5_x0y3, aib4_ch5_x0y3,
                aib3_ch5_x0y3,  aib2_ch5_x0y3,  aib1_ch5_x0y3, aib0_ch5_x0y3,
                aib19_ch5_x0y3, aib18_ch5_x0y3, aib17_ch5_x0y3,aib16_ch5_x0y3,
                aib15_ch5_x0y3, aib14_ch5_x0y3, aib13_ch5_x0y3,aib12_ch5_x0y3,
                aib11_ch5_x0y3, aib10_ch5_x0y3, aib9_ch5_x0y3, aib8_ch5_x0y3,
                aib7_ch5_x0y3,  aib6_ch5_x0y3,  aib5_ch5_x0y3, aib4_ch5_x0y3,
                aib3_ch5_x0y3,  aib2_ch5_x0y3,  aib1_ch5_x0y3, aib0_ch5_x0y3};
*/
    //-----------------------------------------------------------------------------------------
    // Interface instantiation

    dut_io top_io (.i_osc_clk (i_osc_clk), 
                   .i_rx_pma_clk (i_rx_pma_clk),
                   .i_tx_pma_clk (i_tx_pma_clk),
                   .i_cfg_avmm_clk (i_cfg_avmm_clk)
                   );

    //-----------------------------------------------------------------------------------------
    // Testbench instantiation
    test t (top_io);

    aib_top u_aib_top
             (
                    .i_adpt_hard_rst_n           (top_io.i_adpt_hard_rst_n), 
                    .o_rx_xcvrif_rst_n           (),   // FIXME
                    .i_cfg_avmm_clk              (i_cfg_avmm_clk), 
                    .i_cfg_avmm_rst_n            (top_io.i_cfg_avmm_rst_n), 
                    .i_cfg_avmm_addr             (top_io.i_cfg_avmm_addr[16:0]), 
                    .i_cfg_avmm_byte_en          (top_io.i_cfg_avmm_byte_en[3:0]), 
                    .i_cfg_avmm_read             (top_io.i_cfg_avmm_read), 
                    .i_cfg_avmm_write            (top_io.i_cfg_avmm_write), 
                    .i_cfg_avmm_wdata            (top_io.i_cfg_avmm_wdata[31:0]), 
                    .o_cfg_avmm_rdatavld         (o_cfg_avmm_rdatavld),
                    .o_cfg_avmm_rdata            (o_cfg_avmm_rdata), 
                    .o_cfg_avmm_waitreq          (o_cfg_avmm_waitreq), 
                    .i_rx_pma_clk                ({24{i_rx_pma_clk}}), 
                    .i_rx_pma_div2_clk           ({24{i_rx_pma_div2_clk}}), 
                    .i_chnl_ssr                  ({65*24{1'b0}}),   // FIXME
                    .i_rx_pma_data               ({24{top_io.i_rx_pma_data[39:0]}}), 
                    .i_tx_pma_clk                ({24{i_tx_pma_clk}}), 
                    .o_chnl_ssr                  (),        // FIXME 
                    .o_tx_transfer_clk           (o_tx_transfer_clk), 
                    .o_tx_transfer_div2_clk      (o_tx_transfer_div2_clk),        // Not used 
                    .o_tx_pma_data               (o_tx_pma_data_24ch), 
		    .ns_mac_rdy                  ({24{top_io.ns_mac_rdy}}),
                    .ms_sideband                 (ms_sideband),
		    .sl_sideband                 (sl_sideband),
                    .io_aib_ch0                  ({aib95_ch0_x0y0, aib94_ch0_x0y0, 1'b1,          aib94_ch0_x0y0,
                                                   aib91_ch0_x0y0, aib90_ch0_x0y0, aib89_ch0_x0y0,aib88_ch0_x0y0,
                                                   aib87_ch0_x0y0, aib86_ch0_x0y0, aib85_ch0_x0y0,aib84_ch0_x0y0,
                                                   aib85_ch0_x0y0, aib84_ch0_x0y0, aib81_ch0_x0y0,aib80_ch0_x0y0,
                                                   aib79_ch0_x0y0, aib78_ch0_x0y0, aib77_ch0_x0y0,aib76_ch0_x0y0,
                                                   aib75_ch0_x0y0, aib74_ch0_x0y0, aib73_ch0_x0y0,aib72_ch0_x0y0,
                                                   aib71_ch0_x0y0, aib70_ch0_x0y0, aib69_ch0_x0y0,aib68_ch0_x0y0,
                                                   aib67_ch0_x0y0, aib66_ch0_x0y0, 1'b1,          aib64_ch0_x0y0,
                                                   aib63_ch0_x0y0, aib62_ch0_x0y0, 1'b1,          aib60_ch0_x0y0,
                                                   aib59_ch0_x0y0, aib58_ch0_x0y0, aib57_ch0_x0y0,aib56_ch0_x0y0,
                                                   aib55_ch0_x0y0, aib54_ch0_x0y0, aib53_ch0_x0y0,aib52_ch0_x0y0,
                                                   aib51_ch0_x0y0, aib50_ch0_x0y0, aib49_ch0_x0y0,aib48_ch0_x0y0,
                                                   aib47_ch0_x0y0, aib46_ch0_x0y0, aib45_ch0_x0y0,aib44_ch0_x0y0,
                                                   aib41_ch0_x0y0, aib40_ch0_x0y0, aib41_ch0_x0y0,aib40_ch0_x0y0,
                                                   aib19_ch0_x0y0, aib18_ch0_x0y0, aib17_ch0_x0y0,aib16_ch0_x0y0,
                                                   aib15_ch0_x0y0, aib14_ch0_x0y0, aib13_ch0_x0y0,aib12_ch0_x0y0,
                                                   aib11_ch0_x0y0, aib10_ch0_x0y0, aib9_ch0_x0y0, aib8_ch0_x0y0,
                                                   aib7_ch0_x0y0,  aib6_ch0_x0y0,  aib5_ch0_x0y0, aib4_ch0_x0y0,
                                                   aib3_ch0_x0y0,  aib2_ch0_x0y0,  aib1_ch0_x0y0, aib0_ch0_x0y0,
                                                   aib19_ch0_x0y0, aib18_ch0_x0y0, aib17_ch0_x0y0,aib16_ch0_x0y0,
                                                   aib15_ch0_x0y0, aib14_ch0_x0y0, aib13_ch0_x0y0,aib12_ch0_x0y0,
                                                   aib11_ch0_x0y0, aib10_ch0_x0y0, aib9_ch0_x0y0, aib8_ch0_x0y0,
                                                   aib7_ch0_x0y0,  aib6_ch0_x0y0,  aib5_ch0_x0y0, aib4_ch0_x0y0,
                                                   aib3_ch0_x0y0,  aib2_ch0_x0y0,  aib1_ch0_x0y0, aib0_ch0_x0y0}),
                    .io_aib_ch1                  ({aib95_ch1_x0y0, aib94_ch1_x0y0, 1'b1,          aib94_ch1_x0y0,
                                                   aib91_ch1_x0y0, aib90_ch1_x0y0, aib89_ch1_x0y0,aib88_ch1_x0y0,
                                                   aib87_ch1_x0y0, aib86_ch1_x0y0, aib85_ch1_x0y0,aib84_ch1_x0y0,
                                                   aib85_ch1_x0y0, aib84_ch1_x0y0, aib81_ch1_x0y0,aib80_ch1_x0y0,
                                                   aib79_ch1_x0y0, aib78_ch1_x0y0, aib77_ch1_x0y0,aib76_ch1_x0y0,
                                                   aib75_ch1_x0y0, aib74_ch1_x0y0, aib73_ch1_x0y0,aib72_ch1_x0y0,
                                                   aib71_ch1_x0y0, aib70_ch1_x0y0, aib69_ch1_x0y0,aib68_ch1_x0y0,
                                                   aib67_ch1_x0y0, aib66_ch1_x0y0, 1'b1,          aib64_ch1_x0y0,
                                                   aib63_ch1_x0y0, aib62_ch1_x0y0, 1'b1,          aib60_ch1_x0y0,
                                                   aib59_ch1_x0y0, aib58_ch1_x0y0, aib57_ch1_x0y0,aib56_ch1_x0y0,
                                                   aib55_ch1_x0y0, aib54_ch1_x0y0, aib53_ch1_x0y0,aib52_ch1_x0y0,
                                                   aib51_ch1_x0y0, aib50_ch1_x0y0, aib49_ch1_x0y0,aib48_ch1_x0y0,
                                                   aib47_ch1_x0y0, aib46_ch1_x0y0, aib45_ch1_x0y0,aib44_ch1_x0y0,
                                                   aib41_ch1_x0y0, aib40_ch1_x0y0, aib41_ch1_x0y0,aib40_ch1_x0y0,
                                                   aib19_ch1_x0y0, aib18_ch1_x0y0, aib17_ch1_x0y0,aib16_ch1_x0y0,
                                                   aib15_ch1_x0y0, aib14_ch1_x0y0, aib13_ch1_x0y0,aib12_ch1_x0y0,
                                                   aib11_ch1_x0y0, aib10_ch1_x0y0, aib9_ch1_x0y0, aib8_ch1_x0y0,
                                                   aib7_ch1_x0y0,  aib6_ch1_x0y0,  aib5_ch1_x0y0, aib4_ch1_x0y0,
                                                   aib3_ch1_x0y0,  aib2_ch1_x0y0,  aib1_ch1_x0y0, aib0_ch1_x0y0,
                                                   aib19_ch1_x0y0, aib18_ch1_x0y0, aib17_ch1_x0y0,aib16_ch1_x0y0,
                                                   aib15_ch1_x0y0, aib14_ch1_x0y0, aib13_ch1_x0y0,aib12_ch1_x0y0,
                                                   aib11_ch1_x0y0, aib10_ch1_x0y0, aib9_ch1_x0y0, aib8_ch1_x0y0,
                                                   aib7_ch1_x0y0,  aib6_ch1_x0y0,  aib5_ch1_x0y0, aib4_ch1_x0y0,
                                                   aib3_ch1_x0y0,  aib2_ch1_x0y0,  aib1_ch1_x0y0, aib0_ch1_x0y0}),
                    .io_aib_ch2                  ({aib95_ch2_x0y0, aib94_ch2_x0y0, 1'b1,          aib94_ch2_x0y0,
                                                   aib91_ch2_x0y0, aib90_ch2_x0y0, aib89_ch2_x0y0,aib88_ch2_x0y0,
                                                   aib87_ch2_x0y0, aib86_ch2_x0y0, aib85_ch2_x0y0,aib84_ch2_x0y0,
                                                   aib85_ch2_x0y0, aib84_ch2_x0y0, aib81_ch2_x0y0,aib80_ch2_x0y0,
                                                   aib79_ch2_x0y0, aib78_ch2_x0y0, aib77_ch2_x0y0,aib76_ch2_x0y0,
                                                   aib75_ch2_x0y0, aib74_ch2_x0y0, aib73_ch2_x0y0,aib72_ch2_x0y0,
                                                   aib71_ch2_x0y0, aib70_ch2_x0y0, aib69_ch2_x0y0,aib68_ch2_x0y0,
                                                   aib67_ch2_x0y0, aib66_ch2_x0y0, 1'b1,          aib64_ch2_x0y0,
                                                   aib63_ch2_x0y0, aib62_ch2_x0y0, 1'b1,          aib60_ch2_x0y0,
                                                   aib59_ch2_x0y0, aib58_ch2_x0y0, aib57_ch2_x0y0,aib56_ch2_x0y0,
                                                   aib55_ch2_x0y0, aib54_ch2_x0y0, aib53_ch2_x0y0,aib52_ch2_x0y0,
                                                   aib51_ch2_x0y0, aib50_ch2_x0y0, aib49_ch2_x0y0,aib48_ch2_x0y0,
                                                   aib47_ch2_x0y0, aib46_ch2_x0y0, aib45_ch2_x0y0,aib44_ch2_x0y0,
                                                   aib41_ch2_x0y0, aib40_ch2_x0y0, aib41_ch2_x0y0,aib40_ch2_x0y0,
                                                   aib19_ch2_x0y0, aib18_ch2_x0y0, aib17_ch2_x0y0,aib16_ch2_x0y0,
                                                   aib15_ch2_x0y0, aib14_ch2_x0y0, aib13_ch2_x0y0,aib12_ch2_x0y0,
                                                   aib11_ch2_x0y0, aib10_ch2_x0y0, aib9_ch2_x0y0, aib8_ch2_x0y0,
                                                   aib7_ch2_x0y0,  aib6_ch2_x0y0,  aib5_ch2_x0y0, aib4_ch2_x0y0,
                                                   aib3_ch2_x0y0,  aib2_ch2_x0y0,  aib1_ch2_x0y0, aib0_ch2_x0y0,
                                                   aib19_ch2_x0y0, aib18_ch2_x0y0, aib17_ch2_x0y0,aib16_ch2_x0y0,
                                                   aib15_ch2_x0y0, aib14_ch2_x0y0, aib13_ch2_x0y0,aib12_ch2_x0y0,
                                                   aib11_ch2_x0y0, aib10_ch2_x0y0, aib9_ch2_x0y0, aib8_ch2_x0y0,
                                                   aib7_ch2_x0y0,  aib6_ch2_x0y0,  aib5_ch2_x0y0, aib4_ch2_x0y0,
                                                   aib3_ch2_x0y0,  aib2_ch2_x0y0,  aib1_ch2_x0y0, aib0_ch2_x0y0}),
                    .io_aib_ch3                  ({aib95_ch3_x0y0, aib94_ch3_x0y0, 1'b1,          aib94_ch3_x0y0,
                                                   aib91_ch3_x0y0, aib90_ch3_x0y0, aib89_ch3_x0y0,aib88_ch3_x0y0,
                                                   aib87_ch3_x0y0, aib86_ch3_x0y0, aib85_ch3_x0y0,aib84_ch3_x0y0,
                                                   aib85_ch3_x0y0, aib84_ch3_x0y0, aib81_ch3_x0y0,aib80_ch3_x0y0,
                                                   aib79_ch3_x0y0, aib78_ch3_x0y0, aib77_ch3_x0y0,aib76_ch3_x0y0,
                                                   aib75_ch3_x0y0, aib74_ch3_x0y0, aib73_ch3_x0y0,aib72_ch3_x0y0,
                                                   aib71_ch3_x0y0, aib70_ch3_x0y0, aib69_ch3_x0y0,aib68_ch3_x0y0,
                                                   aib67_ch3_x0y0, aib66_ch3_x0y0, 1'b1,          aib64_ch3_x0y0,
                                                   aib63_ch3_x0y0, aib62_ch3_x0y0, 1'b1,          aib60_ch3_x0y0,
                                                   aib59_ch3_x0y0, aib58_ch3_x0y0, aib57_ch3_x0y0,aib56_ch3_x0y0,
                                                   aib55_ch3_x0y0, aib54_ch3_x0y0, aib53_ch3_x0y0,aib52_ch3_x0y0,
                                                   aib51_ch3_x0y0, aib50_ch3_x0y0, aib49_ch3_x0y0,aib48_ch3_x0y0,
                                                   aib47_ch3_x0y0, aib46_ch3_x0y0, aib45_ch3_x0y0,aib44_ch3_x0y0,
                                                   aib41_ch3_x0y0, aib40_ch3_x0y0, aib41_ch3_x0y0,aib40_ch3_x0y0,
                                                   aib19_ch3_x0y0, aib18_ch3_x0y0, aib17_ch3_x0y0,aib16_ch3_x0y0,
                                                   aib15_ch3_x0y0, aib14_ch3_x0y0, aib13_ch3_x0y0,aib12_ch3_x0y0,
                                                   aib11_ch3_x0y0, aib10_ch3_x0y0, aib9_ch3_x0y0, aib8_ch3_x0y0,
                                                   aib7_ch3_x0y0,  aib6_ch3_x0y0,  aib5_ch3_x0y0, aib4_ch3_x0y0,
                                                   aib3_ch3_x0y0,  aib2_ch3_x0y0,  aib1_ch3_x0y0, aib0_ch3_x0y0,
                                                   aib19_ch3_x0y0, aib18_ch3_x0y0, aib17_ch3_x0y0,aib16_ch3_x0y0,
                                                   aib15_ch3_x0y0, aib14_ch3_x0y0, aib13_ch3_x0y0,aib12_ch3_x0y0,
                                                   aib11_ch3_x0y0, aib10_ch3_x0y0, aib9_ch3_x0y0, aib8_ch3_x0y0,
                                                   aib7_ch3_x0y0,  aib6_ch3_x0y0,  aib5_ch3_x0y0, aib4_ch3_x0y0,
                                                   aib3_ch3_x0y0,  aib2_ch3_x0y0,  aib1_ch3_x0y0, aib0_ch3_x0y0}),
                    .io_aib_ch4                  ({aib95_ch4_x0y0, aib94_ch4_x0y0, 1'b1,          aib94_ch4_x0y0,
                                                   aib91_ch4_x0y0, aib90_ch4_x0y0, aib89_ch4_x0y0,aib88_ch4_x0y0,
                                                   aib87_ch4_x0y0, aib86_ch4_x0y0, aib85_ch4_x0y0,aib84_ch4_x0y0,
                                                   aib85_ch4_x0y0, aib84_ch4_x0y0, aib81_ch4_x0y0,aib80_ch4_x0y0,
                                                   aib79_ch4_x0y0, aib78_ch4_x0y0, aib77_ch4_x0y0,aib76_ch4_x0y0,
                                                   aib75_ch4_x0y0, aib74_ch4_x0y0, aib73_ch4_x0y0,aib72_ch4_x0y0,
                                                   aib71_ch4_x0y0, aib70_ch4_x0y0, aib69_ch4_x0y0,aib68_ch4_x0y0,
                                                   aib67_ch4_x0y0, aib66_ch4_x0y0, 1'b1,          aib64_ch4_x0y0,
                                                   aib63_ch4_x0y0, aib62_ch4_x0y0, 1'b1,          aib60_ch4_x0y0,
                                                   aib59_ch4_x0y0, aib58_ch4_x0y0, aib57_ch4_x0y0,aib56_ch4_x0y0,
                                                   aib55_ch4_x0y0, aib54_ch4_x0y0, aib53_ch4_x0y0,aib52_ch4_x0y0,
                                                   aib51_ch4_x0y0, aib50_ch4_x0y0, aib49_ch4_x0y0,aib48_ch4_x0y0,
                                                   aib47_ch4_x0y0, aib46_ch4_x0y0, aib45_ch4_x0y0,aib44_ch4_x0y0,
                                                   aib41_ch4_x0y0, aib40_ch4_x0y0, aib41_ch4_x0y0,aib40_ch4_x0y0,
                                                   aib19_ch4_x0y0, aib18_ch4_x0y0, aib17_ch4_x0y0,aib16_ch4_x0y0,
                                                   aib15_ch4_x0y0, aib14_ch4_x0y0, aib13_ch4_x0y0,aib12_ch4_x0y0,
                                                   aib11_ch4_x0y0, aib10_ch4_x0y0, aib9_ch4_x0y0, aib8_ch4_x0y0,
                                                   aib7_ch4_x0y0,  aib6_ch4_x0y0,  aib5_ch4_x0y0, aib4_ch4_x0y0,
                                                   aib3_ch4_x0y0,  aib2_ch4_x0y0,  aib1_ch4_x0y0, aib0_ch4_x0y0,
                                                   aib19_ch4_x0y0, aib18_ch4_x0y0, aib17_ch4_x0y0,aib16_ch4_x0y0,
                                                   aib15_ch4_x0y0, aib14_ch4_x0y0, aib13_ch4_x0y0,aib12_ch4_x0y0,
                                                   aib11_ch4_x0y0, aib10_ch4_x0y0, aib9_ch4_x0y0, aib8_ch4_x0y0,
                                                   aib7_ch4_x0y0,  aib6_ch4_x0y0,  aib5_ch4_x0y0, aib4_ch4_x0y0,
                                                   aib3_ch4_x0y0,  aib2_ch4_x0y0,  aib1_ch4_x0y0, aib0_ch4_x0y0}),
                    .io_aib_ch5                  ({aib95_ch5_x0y0, aib94_ch5_x0y0, 1'b1,          aib94_ch5_x0y0,
                                                   aib91_ch5_x0y0, aib90_ch5_x0y0, aib89_ch5_x0y0,aib88_ch5_x0y0,
                                                   aib87_ch5_x0y0, aib86_ch5_x0y0, aib85_ch5_x0y0,aib84_ch5_x0y0,
                                                   aib85_ch5_x0y0, aib84_ch5_x0y0, aib81_ch5_x0y0,aib80_ch5_x0y0,
                                                   aib79_ch5_x0y0, aib78_ch5_x0y0, aib77_ch5_x0y0,aib76_ch5_x0y0,
                                                   aib75_ch5_x0y0, aib74_ch5_x0y0, aib73_ch5_x0y0,aib72_ch5_x0y0,
                                                   aib71_ch5_x0y0, aib70_ch5_x0y0, aib69_ch5_x0y0,aib68_ch5_x0y0,
                                                   aib67_ch5_x0y0, aib66_ch5_x0y0, 1'b1,          aib64_ch5_x0y0,
                                                   aib63_ch5_x0y0, aib62_ch5_x0y0, 1'b1,          aib60_ch5_x0y0,
                                                   aib59_ch5_x0y0, aib58_ch5_x0y0, aib57_ch5_x0y0,aib56_ch5_x0y0,
                                                   aib55_ch5_x0y0, aib54_ch5_x0y0, aib53_ch5_x0y0,aib52_ch5_x0y0,
                                                   aib51_ch5_x0y0, aib50_ch5_x0y0, aib49_ch5_x0y0,aib48_ch5_x0y0,
                                                   aib47_ch5_x0y0, aib46_ch5_x0y0, aib45_ch5_x0y0,aib44_ch5_x0y0,
                                                   aib41_ch5_x0y0, aib40_ch5_x0y0, aib41_ch5_x0y0,aib40_ch5_x0y0,
                                                   aib19_ch5_x0y0, aib18_ch5_x0y0, aib17_ch5_x0y0,aib16_ch5_x0y0,
                                                   aib15_ch5_x0y0, aib14_ch5_x0y0, aib13_ch5_x0y0,aib12_ch5_x0y0,
                                                   aib11_ch5_x0y0, aib10_ch5_x0y0, aib9_ch5_x0y0, aib8_ch5_x0y0,
                                                   aib7_ch5_x0y0,  aib6_ch5_x0y0,  aib5_ch5_x0y0, aib4_ch5_x0y0,
                                                   aib3_ch5_x0y0,  aib2_ch5_x0y0,  aib1_ch5_x0y0, aib0_ch5_x0y0,
                                                   aib19_ch5_x0y0, aib18_ch5_x0y0, aib17_ch5_x0y0,aib16_ch5_x0y0,
                                                   aib15_ch5_x0y0, aib14_ch5_x0y0, aib13_ch5_x0y0,aib12_ch5_x0y0,
                                                   aib11_ch5_x0y0, aib10_ch5_x0y0, aib9_ch5_x0y0, aib8_ch5_x0y0,
                                                   aib7_ch5_x0y0,  aib6_ch5_x0y0,  aib5_ch5_x0y0, aib4_ch5_x0y0,
                                                   aib3_ch5_x0y0,  aib2_ch5_x0y0,  aib1_ch5_x0y0, aib0_ch5_x0y0}),
                    .io_aib_ch6                  ({aib95_ch0_x0y1, aib94_ch0_x0y1, 1'b1,          aib94_ch0_x0y1,
                                                   aib91_ch0_x0y1, aib90_ch0_x0y1, aib89_ch0_x0y1,aib88_ch0_x0y1,
                                                   aib87_ch0_x0y1, aib86_ch0_x0y1, aib85_ch0_x0y1,aib84_ch0_x0y1,
                                                   aib85_ch0_x0y1, aib84_ch0_x0y1, aib81_ch0_x0y1,aib80_ch0_x0y1,
                                                   aib79_ch0_x0y1, aib78_ch0_x0y1, aib77_ch0_x0y1,aib76_ch0_x0y1,
                                                   aib75_ch0_x0y1, aib74_ch0_x0y1, aib73_ch0_x0y1,aib72_ch0_x0y1,
                                                   aib71_ch0_x0y1, aib70_ch0_x0y1, aib69_ch0_x0y1,aib68_ch0_x0y1,
                                                   aib67_ch0_x0y1, aib66_ch0_x0y1, 1'b1,          aib64_ch0_x0y1,
                                                   aib63_ch0_x0y1, aib62_ch0_x0y1, 1'b1,          aib60_ch0_x0y1,
                                                   aib59_ch0_x0y1, aib58_ch0_x0y1, aib57_ch0_x0y1,aib56_ch0_x0y1,
                                                   aib55_ch0_x0y1, aib54_ch0_x0y1, aib53_ch0_x0y1,aib52_ch0_x0y1,
                                                   aib51_ch0_x0y1, aib50_ch0_x0y1, aib49_ch0_x0y1,aib48_ch0_x0y1,
                                                   aib47_ch0_x0y1, aib46_ch0_x0y1, aib45_ch0_x0y1,aib44_ch0_x0y1,
                                                   aib41_ch0_x0y1, aib40_ch0_x0y1, aib41_ch0_x0y1,aib40_ch0_x0y1,
                                                   aib19_ch0_x0y1, aib18_ch0_x0y1, aib17_ch0_x0y1,aib16_ch0_x0y1,
                                                   aib15_ch0_x0y1, aib14_ch0_x0y1, aib13_ch0_x0y1,aib12_ch0_x0y1,
                                                   aib11_ch0_x0y1, aib10_ch0_x0y1, aib9_ch0_x0y1, aib8_ch0_x0y1,
                                                   aib7_ch0_x0y1,  aib6_ch0_x0y1,  aib5_ch0_x0y1, aib4_ch0_x0y1,
                                                   aib3_ch0_x0y1,  aib2_ch0_x0y1,  aib1_ch0_x0y1, aib0_ch0_x0y1,
                                                   aib19_ch0_x0y1, aib18_ch0_x0y1, aib17_ch0_x0y1,aib16_ch0_x0y1,
                                                   aib15_ch0_x0y1, aib14_ch0_x0y1, aib13_ch0_x0y1,aib12_ch0_x0y1,
                                                   aib11_ch0_x0y1, aib10_ch0_x0y1, aib9_ch0_x0y1, aib8_ch0_x0y1,
                                                   aib7_ch0_x0y1,  aib6_ch0_x0y1,  aib5_ch0_x0y1, aib4_ch0_x0y1,
                                                   aib3_ch0_x0y1,  aib2_ch0_x0y1,  aib1_ch0_x0y1, aib0_ch0_x0y1}),
                    .io_aib_ch7                  ({aib95_ch1_x0y1, aib94_ch1_x0y1, 1'b1,          aib94_ch1_x0y1,
                                                   aib91_ch1_x0y1, aib90_ch1_x0y1, aib89_ch1_x0y1,aib88_ch1_x0y1,
                                                   aib87_ch1_x0y1, aib86_ch1_x0y1, aib85_ch1_x0y1,aib84_ch1_x0y1,
                                                   aib85_ch1_x0y1, aib84_ch1_x0y1, aib81_ch1_x0y1,aib80_ch1_x0y1,
                                                   aib79_ch1_x0y1, aib78_ch1_x0y1, aib77_ch1_x0y1,aib76_ch1_x0y1,
                                                   aib75_ch1_x0y1, aib74_ch1_x0y1, aib73_ch1_x0y1,aib72_ch1_x0y1,
                                                   aib71_ch1_x0y1, aib70_ch1_x0y1, aib69_ch1_x0y1,aib68_ch1_x0y1,
                                                   aib67_ch1_x0y1, aib66_ch1_x0y1, 1'b1,          aib64_ch1_x0y1,
                                                   aib63_ch1_x0y1, aib62_ch1_x0y1, 1'b1,          aib60_ch1_x0y1,
                                                   aib59_ch1_x0y1, aib58_ch1_x0y1, aib57_ch1_x0y1,aib56_ch1_x0y1,
                                                   aib55_ch1_x0y1, aib54_ch1_x0y1, aib53_ch1_x0y1,aib52_ch1_x0y1,
                                                   aib51_ch1_x0y1, aib50_ch1_x0y1, aib49_ch1_x0y1,aib48_ch1_x0y1,
                                                   aib47_ch1_x0y1, aib46_ch1_x0y1, aib45_ch1_x0y1,aib44_ch1_x0y1,
                                                   aib41_ch1_x0y1, aib40_ch1_x0y1, aib41_ch1_x0y1,aib40_ch1_x0y1,
                                                   aib19_ch1_x0y1, aib18_ch1_x0y1, aib17_ch1_x0y1,aib16_ch1_x0y1,
                                                   aib15_ch1_x0y1, aib14_ch1_x0y1, aib13_ch1_x0y1,aib12_ch1_x0y1,
                                                   aib11_ch1_x0y1, aib10_ch1_x0y1, aib9_ch1_x0y1, aib8_ch1_x0y1,
                                                   aib7_ch1_x0y1,  aib6_ch1_x0y1,  aib5_ch1_x0y1, aib4_ch1_x0y1,
                                                   aib3_ch1_x0y1,  aib2_ch1_x0y1,  aib1_ch1_x0y1, aib0_ch1_x0y1,
                                                   aib19_ch1_x0y1, aib18_ch1_x0y1, aib17_ch1_x0y1,aib16_ch1_x0y1,
                                                   aib15_ch1_x0y1, aib14_ch1_x0y1, aib13_ch1_x0y1,aib12_ch1_x0y1,
                                                   aib11_ch1_x0y1, aib10_ch1_x0y1, aib9_ch1_x0y1, aib8_ch1_x0y1,
                                                   aib7_ch1_x0y1,  aib6_ch1_x0y1,  aib5_ch1_x0y1, aib4_ch1_x0y1,
                                                   aib3_ch1_x0y1,  aib2_ch1_x0y1,  aib1_ch1_x0y1, aib0_ch1_x0y1}),
                    .io_aib_ch8                  ({aib95_ch2_x0y1, aib94_ch2_x0y1, 1'b1,          aib94_ch2_x0y1,
                                                   aib91_ch2_x0y1, aib90_ch2_x0y1, aib89_ch2_x0y1,aib88_ch2_x0y1,
                                                   aib87_ch2_x0y1, aib86_ch2_x0y1, aib85_ch2_x0y1,aib84_ch2_x0y1,
                                                   aib85_ch2_x0y1, aib84_ch2_x0y1, aib81_ch2_x0y1,aib80_ch2_x0y1,
                                                   aib79_ch2_x0y1, aib78_ch2_x0y1, aib77_ch2_x0y1,aib76_ch2_x0y1,
                                                   aib75_ch2_x0y1, aib74_ch2_x0y1, aib73_ch2_x0y1,aib72_ch2_x0y1,
                                                   aib71_ch2_x0y1, aib70_ch2_x0y1, aib69_ch2_x0y1,aib68_ch2_x0y1,
                                                   aib67_ch2_x0y1, aib66_ch2_x0y1, 1'b1,          aib64_ch2_x0y1,
                                                   aib63_ch2_x0y1, aib62_ch2_x0y1, 1'b1,          aib60_ch2_x0y1,
                                                   aib59_ch2_x0y1, aib58_ch2_x0y1, aib57_ch2_x0y1,aib56_ch2_x0y1,
                                                   aib55_ch2_x0y1, aib54_ch2_x0y1, aib53_ch2_x0y1,aib52_ch2_x0y1,
                                                   aib51_ch2_x0y1, aib50_ch2_x0y1, aib49_ch2_x0y1,aib48_ch2_x0y1,
                                                   aib47_ch2_x0y1, aib46_ch2_x0y1, aib45_ch2_x0y1,aib44_ch2_x0y1,
                                                   aib41_ch2_x0y1, aib40_ch2_x0y1, aib41_ch2_x0y1,aib40_ch2_x0y1,
                                                   aib19_ch2_x0y1, aib18_ch2_x0y1, aib17_ch2_x0y1,aib16_ch2_x0y1,
                                                   aib15_ch2_x0y1, aib14_ch2_x0y1, aib13_ch2_x0y1,aib12_ch2_x0y1,
                                                   aib11_ch2_x0y1, aib10_ch2_x0y1, aib9_ch2_x0y1, aib8_ch2_x0y1,
                                                   aib7_ch2_x0y1,  aib6_ch2_x0y1,  aib5_ch2_x0y1, aib4_ch2_x0y1,
                                                   aib3_ch2_x0y1,  aib2_ch2_x0y1,  aib1_ch2_x0y1, aib0_ch2_x0y1,
                                                   aib19_ch2_x0y1, aib18_ch2_x0y1, aib17_ch2_x0y1,aib16_ch2_x0y1,
                                                   aib15_ch2_x0y1, aib14_ch2_x0y1, aib13_ch2_x0y1,aib12_ch2_x0y1,
                                                   aib11_ch2_x0y1, aib10_ch2_x0y1, aib9_ch2_x0y1, aib8_ch2_x0y1,
                                                   aib7_ch2_x0y1,  aib6_ch2_x0y1,  aib5_ch2_x0y1, aib4_ch2_x0y1,
                                                   aib3_ch2_x0y1,  aib2_ch2_x0y1,  aib1_ch2_x0y1, aib0_ch2_x0y1}),
                    .io_aib_ch9                  ({aib95_ch3_x0y1, aib94_ch3_x0y1, 1'b1,          aib94_ch3_x0y1,
                                                   aib91_ch3_x0y1, aib90_ch3_x0y1, aib89_ch3_x0y1,aib88_ch3_x0y1,
                                                   aib87_ch3_x0y1, aib86_ch3_x0y1, aib85_ch3_x0y1,aib84_ch3_x0y1,
                                                   aib85_ch3_x0y1, aib84_ch3_x0y1, aib81_ch3_x0y1,aib80_ch3_x0y1,
                                                   aib79_ch3_x0y1, aib78_ch3_x0y1, aib77_ch3_x0y1,aib76_ch3_x0y1,
                                                   aib75_ch3_x0y1, aib74_ch3_x0y1, aib73_ch3_x0y1,aib72_ch3_x0y1,
                                                   aib71_ch3_x0y1, aib70_ch3_x0y1, aib69_ch3_x0y1,aib68_ch3_x0y1,
                                                   aib67_ch3_x0y1, aib66_ch3_x0y1, 1'b1,          aib64_ch3_x0y1,
                                                   aib63_ch3_x0y1, aib62_ch3_x0y1, 1'b1,          aib60_ch3_x0y1,
                                                   aib59_ch3_x0y1, aib58_ch3_x0y1, aib57_ch3_x0y1,aib56_ch3_x0y1,
                                                   aib55_ch3_x0y1, aib54_ch3_x0y1, aib53_ch3_x0y1,aib52_ch3_x0y1,
                                                   aib51_ch3_x0y1, aib50_ch3_x0y1, aib49_ch3_x0y1,aib48_ch3_x0y1,
                                                   aib47_ch3_x0y1, aib46_ch3_x0y1, aib45_ch3_x0y1,aib44_ch3_x0y1,
                                                   aib41_ch3_x0y1, aib40_ch3_x0y1, aib41_ch3_x0y1,aib40_ch3_x0y1,
                                                   aib19_ch3_x0y1, aib18_ch3_x0y1, aib17_ch3_x0y1,aib16_ch3_x0y1,
                                                   aib15_ch3_x0y1, aib14_ch3_x0y1, aib13_ch3_x0y1,aib12_ch3_x0y1,
                                                   aib11_ch3_x0y1, aib10_ch3_x0y1, aib9_ch3_x0y1, aib8_ch3_x0y1,
                                                   aib7_ch3_x0y1,  aib6_ch3_x0y1,  aib5_ch3_x0y1, aib4_ch3_x0y1,
                                                   aib3_ch3_x0y1,  aib2_ch3_x0y1,  aib1_ch3_x0y1, aib0_ch3_x0y1,
                                                   aib19_ch3_x0y1, aib18_ch3_x0y1, aib17_ch3_x0y1,aib16_ch3_x0y1,
                                                   aib15_ch3_x0y1, aib14_ch3_x0y1, aib13_ch3_x0y1,aib12_ch3_x0y1,
                                                   aib11_ch3_x0y1, aib10_ch3_x0y1, aib9_ch3_x0y1, aib8_ch3_x0y1,
                                                   aib7_ch3_x0y1,  aib6_ch3_x0y1,  aib5_ch3_x0y1, aib4_ch3_x0y1,
                                                   aib3_ch3_x0y1,  aib2_ch3_x0y1,  aib1_ch3_x0y1, aib0_ch3_x0y1}),
                    .io_aib_ch10                 ({aib95_ch4_x0y1, aib94_ch4_x0y1, 1'b1,         aib94_ch4_x0y1,
                                                   aib91_ch4_x0y1, aib90_ch4_x0y1, aib89_ch4_x0y1,aib88_ch4_x0y1,
                                                   aib87_ch4_x0y1, aib86_ch4_x0y1, aib85_ch4_x0y1,aib84_ch4_x0y1,
                                                   aib85_ch4_x0y1, aib84_ch4_x0y1, aib81_ch4_x0y1,aib80_ch4_x0y1,
                                                   aib79_ch4_x0y1, aib78_ch4_x0y1, aib77_ch4_x0y1,aib76_ch4_x0y1,
                                                   aib75_ch4_x0y1, aib74_ch4_x0y1, aib73_ch4_x0y1,aib72_ch4_x0y1,
                                                   aib71_ch4_x0y1, aib70_ch4_x0y1, aib69_ch4_x0y1,aib68_ch4_x0y1,
                                                   aib67_ch4_x0y1, aib66_ch4_x0y1, 1'b1,          aib64_ch4_x0y1,
                                                   aib63_ch4_x0y1, aib62_ch4_x0y1, 1'b1,          aib60_ch4_x0y1,
                                                   aib59_ch4_x0y1, aib58_ch4_x0y1, aib57_ch4_x0y1,aib56_ch4_x0y1,
                                                   aib55_ch4_x0y1, aib54_ch4_x0y1, aib53_ch4_x0y1,aib52_ch4_x0y1,
                                                   aib51_ch4_x0y1, aib50_ch4_x0y1, aib49_ch4_x0y1,aib48_ch4_x0y1,
                                                   aib47_ch4_x0y1, aib46_ch4_x0y1, aib45_ch4_x0y1,aib44_ch4_x0y1,
                                                   aib41_ch4_x0y1, aib40_ch4_x0y1, aib41_ch4_x0y1,aib40_ch4_x0y1,
                                                   aib19_ch4_x0y1, aib18_ch4_x0y1, aib17_ch4_x0y1,aib16_ch4_x0y1,
                                                   aib15_ch4_x0y1, aib14_ch4_x0y1, aib13_ch4_x0y1,aib12_ch4_x0y1,
                                                   aib11_ch4_x0y1, aib10_ch4_x0y1, aib9_ch4_x0y1, aib8_ch4_x0y1,
                                                   aib7_ch4_x0y1,  aib6_ch4_x0y1,  aib5_ch4_x0y1, aib4_ch4_x0y1,
                                                   aib3_ch4_x0y1,  aib2_ch4_x0y1,  aib1_ch4_x0y1, aib0_ch4_x0y1,
                                                   aib19_ch4_x0y1, aib18_ch4_x0y1, aib17_ch4_x0y1,aib16_ch4_x0y1,
                                                   aib15_ch4_x0y1, aib14_ch4_x0y1, aib13_ch4_x0y1,aib12_ch4_x0y1,
                                                   aib11_ch4_x0y1, aib10_ch4_x0y1, aib9_ch4_x0y1, aib8_ch4_x0y1,
                                                   aib7_ch4_x0y1,  aib6_ch4_x0y1,  aib5_ch4_x0y1, aib4_ch4_x0y1,
                                                   aib3_ch4_x0y1,  aib2_ch4_x0y1,  aib1_ch4_x0y1, aib0_ch4_x0y1}),
                    .io_aib_ch11                 ({aib95_ch5_x0y1, aib94_ch5_x0y1, 1'b1,         aib94_ch5_x0y1,
                                                   aib91_ch5_x0y1, aib90_ch5_x0y1, aib89_ch5_x0y1,aib88_ch5_x0y1,
                                                   aib87_ch5_x0y1, aib86_ch5_x0y1, aib85_ch5_x0y1,aib84_ch5_x0y1,
                                                   aib85_ch5_x0y1, aib84_ch5_x0y1, aib81_ch5_x0y1,aib80_ch5_x0y1,
                                                   aib79_ch5_x0y1, aib78_ch5_x0y1, aib77_ch5_x0y1,aib76_ch5_x0y1,
                                                   aib75_ch5_x0y1, aib74_ch5_x0y1, aib73_ch5_x0y1,aib72_ch5_x0y1,
                                                   aib71_ch5_x0y1, aib70_ch5_x0y1, aib69_ch5_x0y1,aib68_ch5_x0y1,
                                                   aib67_ch5_x0y1, aib66_ch5_x0y1, 1'b1,          aib64_ch5_x0y1,
                                                   aib63_ch5_x0y1, aib62_ch5_x0y1, 1'b1,          aib60_ch5_x0y1,
                                                   aib59_ch5_x0y1, aib58_ch5_x0y1, aib57_ch5_x0y1,aib56_ch5_x0y1,
                                                   aib55_ch5_x0y1, aib54_ch5_x0y1, aib53_ch5_x0y1,aib52_ch5_x0y1,
                                                   aib51_ch5_x0y1, aib50_ch5_x0y1, aib49_ch5_x0y1,aib48_ch5_x0y1,
                                                   aib47_ch5_x0y1, aib46_ch5_x0y1, aib45_ch5_x0y1,aib44_ch5_x0y1,
                                                   aib41_ch5_x0y1, aib40_ch5_x0y1, aib41_ch5_x0y1,aib40_ch5_x0y1,
                                                   aib19_ch5_x0y1, aib18_ch5_x0y1, aib17_ch5_x0y1,aib16_ch5_x0y1,
                                                   aib15_ch5_x0y1, aib14_ch5_x0y1, aib13_ch5_x0y1,aib12_ch5_x0y1,
                                                   aib11_ch5_x0y1, aib10_ch5_x0y1, aib9_ch5_x0y1, aib8_ch5_x0y1,
                                                   aib7_ch5_x0y1,  aib6_ch5_x0y1,  aib5_ch5_x0y1, aib4_ch5_x0y1,
                                                   aib3_ch5_x0y1,  aib2_ch5_x0y1,  aib1_ch5_x0y1, aib0_ch5_x0y1,
                                                   aib19_ch5_x0y1, aib18_ch5_x0y1, aib17_ch5_x0y1,aib16_ch5_x0y1,
                                                   aib15_ch5_x0y1, aib14_ch5_x0y1, aib13_ch5_x0y1,aib12_ch5_x0y1,
                                                   aib11_ch5_x0y1, aib10_ch5_x0y1, aib9_ch5_x0y1, aib8_ch5_x0y1,
                                                   aib7_ch5_x0y1,  aib6_ch5_x0y1,  aib5_ch5_x0y1, aib4_ch5_x0y1,
                                                   aib3_ch5_x0y1,  aib2_ch5_x0y1,  aib1_ch5_x0y1, aib0_ch5_x0y1}),
                    .io_aib_ch12                 ({aib95_ch0_x0y2, aib94_ch0_x0y2, 1'b1,         aib94_ch0_x0y2,
                                                   aib91_ch0_x0y2, aib90_ch0_x0y2, aib89_ch0_x0y2,aib88_ch0_x0y2,
                                                   aib87_ch0_x0y2, aib86_ch0_x0y2, aib85_ch0_x0y2,aib84_ch0_x0y2,
                                                   aib85_ch0_x0y2, aib84_ch0_x0y2, aib81_ch0_x0y2,aib80_ch0_x0y2,
                                                   aib79_ch0_x0y2, aib78_ch0_x0y2, aib77_ch0_x0y2,aib76_ch0_x0y2,
                                                   aib75_ch0_x0y2, aib74_ch0_x0y2, aib73_ch0_x0y2,aib72_ch0_x0y2,
                                                   aib71_ch0_x0y2, aib70_ch0_x0y2, aib69_ch0_x0y2,aib68_ch0_x0y2,
                                                   aib67_ch0_x0y2, aib66_ch0_x0y2, 1'b1,          aib64_ch0_x0y2,
                                                   aib63_ch0_x0y2, aib62_ch0_x0y2, 1'b1,          aib60_ch0_x0y2,
                                                   aib59_ch0_x0y2, aib58_ch0_x0y2, aib57_ch0_x0y2,aib56_ch0_x0y2,
                                                   aib55_ch0_x0y2, aib54_ch0_x0y2, aib53_ch0_x0y2,aib52_ch0_x0y2,
                                                   aib51_ch0_x0y2, aib50_ch0_x0y2, aib49_ch0_x0y2,aib48_ch0_x0y2,
                                                   aib47_ch0_x0y2, aib46_ch0_x0y2, aib45_ch0_x0y2,aib44_ch0_x0y2,
                                                   aib41_ch0_x0y2, aib40_ch0_x0y2, aib41_ch0_x0y2,aib40_ch0_x0y2,
                                                   aib19_ch0_x0y2, aib18_ch0_x0y2, aib17_ch0_x0y2,aib16_ch0_x0y2,
                                                   aib15_ch0_x0y2, aib14_ch0_x0y2, aib13_ch0_x0y2,aib12_ch0_x0y2,
                                                   aib11_ch0_x0y2, aib10_ch0_x0y2, aib9_ch0_x0y2, aib8_ch0_x0y2,
                                                   aib7_ch0_x0y2,  aib6_ch0_x0y2,  aib5_ch0_x0y2, aib4_ch0_x0y2,
                                                   aib3_ch0_x0y2,  aib2_ch0_x0y2,  aib1_ch0_x0y2, aib0_ch0_x0y2,
                                                   aib19_ch0_x0y2, aib18_ch0_x0y2, aib17_ch0_x0y2,aib16_ch0_x0y2,
                                                   aib15_ch0_x0y2, aib14_ch0_x0y2, aib13_ch0_x0y2,aib12_ch0_x0y2,
                                                   aib11_ch0_x0y2, aib10_ch0_x0y2, aib9_ch0_x0y2, aib8_ch0_x0y2,
                                                   aib7_ch0_x0y2,  aib6_ch0_x0y2,  aib5_ch0_x0y2, aib4_ch0_x0y2,
                                                   aib3_ch0_x0y2,  aib2_ch0_x0y2,  aib1_ch0_x0y2, aib0_ch0_x0y2}),
                    .io_aib_ch13                 ({aib95_ch1_x0y2, aib94_ch1_x0y2, 1'b1,         aib94_ch1_x0y2,
                                                   aib91_ch1_x0y2, aib90_ch1_x0y2, aib89_ch1_x0y2,aib88_ch1_x0y2,
                                                   aib87_ch1_x0y2, aib86_ch1_x0y2, aib85_ch1_x0y2,aib84_ch1_x0y2,
                                                   aib85_ch1_x0y2, aib84_ch1_x0y2, aib81_ch1_x0y2,aib80_ch1_x0y2,
                                                   aib79_ch1_x0y2, aib78_ch1_x0y2, aib77_ch1_x0y2,aib76_ch1_x0y2,
                                                   aib75_ch1_x0y2, aib74_ch1_x0y2, aib73_ch1_x0y2,aib72_ch1_x0y2,
                                                   aib71_ch1_x0y2, aib70_ch1_x0y2, aib69_ch1_x0y2,aib68_ch1_x0y2,
                                                   aib67_ch1_x0y2, aib66_ch1_x0y2, 1'b1,          aib64_ch1_x0y2,
                                                   aib63_ch1_x0y2, aib62_ch1_x0y2, 1'b1,          aib60_ch1_x0y2,
                                                   aib59_ch1_x0y2, aib58_ch1_x0y2, aib57_ch1_x0y2,aib56_ch1_x0y2,
                                                   aib55_ch1_x0y2, aib54_ch1_x0y2, aib53_ch1_x0y2,aib52_ch1_x0y2,
                                                   aib51_ch1_x0y2, aib50_ch1_x0y2, aib49_ch1_x0y2,aib48_ch1_x0y2,
                                                   aib47_ch1_x0y2, aib46_ch1_x0y2, aib45_ch1_x0y2,aib44_ch1_x0y2,
                                                   aib41_ch1_x0y2, aib40_ch1_x0y2, aib41_ch1_x0y2,aib40_ch1_x0y2,
                                                   aib19_ch1_x0y2, aib18_ch1_x0y2, aib17_ch1_x0y2,aib16_ch1_x0y2,
                                                   aib15_ch1_x0y2, aib14_ch1_x0y2, aib13_ch1_x0y2,aib12_ch1_x0y2,
                                                   aib11_ch1_x0y2, aib10_ch1_x0y2, aib9_ch1_x0y2, aib8_ch1_x0y2,
                                                   aib7_ch1_x0y2,  aib6_ch1_x0y2,  aib5_ch1_x0y2, aib4_ch1_x0y2,
                                                   aib3_ch1_x0y2,  aib2_ch1_x0y2,  aib1_ch1_x0y2, aib0_ch1_x0y2,
                                                   aib19_ch1_x0y2, aib18_ch1_x0y2, aib17_ch1_x0y2,aib16_ch1_x0y2,
                                                   aib15_ch1_x0y2, aib14_ch1_x0y2, aib13_ch1_x0y2,aib12_ch1_x0y2,
                                                   aib11_ch1_x0y2, aib10_ch1_x0y2, aib9_ch1_x0y2, aib8_ch1_x0y2,
                                                   aib7_ch1_x0y2,  aib6_ch1_x0y2,  aib5_ch1_x0y2, aib4_ch1_x0y2,
                                                   aib3_ch1_x0y2,  aib2_ch1_x0y2,  aib1_ch1_x0y2, aib0_ch1_x0y2}),
                    .io_aib_ch14                 ({aib95_ch2_x0y2, aib94_ch2_x0y2, 1'b1,         aib94_ch2_x0y2,
                                                   aib91_ch2_x0y2, aib90_ch2_x0y2, aib89_ch2_x0y2,aib88_ch2_x0y2,
                                                   aib87_ch2_x0y2, aib86_ch2_x0y2, aib85_ch2_x0y2,aib84_ch2_x0y2,
                                                   aib85_ch2_x0y2, aib84_ch2_x0y2, aib81_ch2_x0y2,aib80_ch2_x0y2,
                                                   aib79_ch2_x0y2, aib78_ch2_x0y2, aib77_ch2_x0y2,aib76_ch2_x0y2,
                                                   aib75_ch2_x0y2, aib74_ch2_x0y2, aib73_ch2_x0y2,aib72_ch2_x0y2,
                                                   aib71_ch2_x0y2, aib70_ch2_x0y2, aib69_ch2_x0y2,aib68_ch2_x0y2,
                                                   aib67_ch2_x0y2, aib66_ch2_x0y2, 1'b1,          aib64_ch2_x0y2,
                                                   aib63_ch2_x0y2, aib62_ch2_x0y2, 1'b1,          aib60_ch2_x0y2,
                                                   aib59_ch2_x0y2, aib58_ch2_x0y2, aib57_ch2_x0y2,aib56_ch2_x0y2,
                                                   aib55_ch2_x0y2, aib54_ch2_x0y2, aib53_ch2_x0y2,aib52_ch2_x0y2,
                                                   aib51_ch2_x0y2, aib50_ch2_x0y2, aib49_ch2_x0y2,aib48_ch2_x0y2,
                                                   aib47_ch2_x0y2, aib46_ch2_x0y2, aib45_ch2_x0y2,aib44_ch2_x0y2,
                                                   aib41_ch2_x0y2, aib40_ch2_x0y2, aib41_ch2_x0y2,aib40_ch2_x0y2,
                                                   aib19_ch2_x0y2, aib18_ch2_x0y2, aib17_ch2_x0y2,aib16_ch2_x0y2,
                                                   aib15_ch2_x0y2, aib14_ch2_x0y2, aib13_ch2_x0y2,aib12_ch2_x0y2,
                                                   aib11_ch2_x0y2, aib10_ch2_x0y2, aib9_ch2_x0y2, aib8_ch2_x0y2,
                                                   aib7_ch2_x0y2,  aib6_ch2_x0y2,  aib5_ch2_x0y2, aib4_ch2_x0y2,
                                                   aib3_ch2_x0y2,  aib2_ch2_x0y2,  aib1_ch2_x0y2, aib0_ch2_x0y2,
                                                   aib19_ch2_x0y2, aib18_ch2_x0y2, aib17_ch2_x0y2,aib16_ch2_x0y2,
                                                   aib15_ch2_x0y2, aib14_ch2_x0y2, aib13_ch2_x0y2,aib12_ch2_x0y2,
                                                   aib11_ch2_x0y2, aib10_ch2_x0y2, aib9_ch2_x0y2, aib8_ch2_x0y2,
                                                   aib7_ch2_x0y2,  aib6_ch2_x0y2,  aib5_ch2_x0y2, aib4_ch2_x0y2,
                                                   aib3_ch2_x0y2,  aib2_ch2_x0y2,  aib1_ch2_x0y2, aib0_ch2_x0y2}),
                    .io_aib_ch15                 ({aib95_ch3_x0y2, aib94_ch3_x0y2, 1'b1,         aib94_ch3_x0y2,
                                                   aib91_ch3_x0y2, aib90_ch3_x0y2, aib89_ch3_x0y2,aib88_ch3_x0y2,
                                                   aib87_ch3_x0y2, aib86_ch3_x0y2, aib85_ch3_x0y2,aib84_ch3_x0y2,
                                                   aib85_ch3_x0y2, aib84_ch3_x0y2, aib81_ch3_x0y2,aib80_ch3_x0y2,
                                                   aib79_ch3_x0y2, aib78_ch3_x0y2, aib77_ch3_x0y2,aib76_ch3_x0y2,
                                                   aib75_ch3_x0y2, aib74_ch3_x0y2, aib73_ch3_x0y2,aib72_ch3_x0y2,
                                                   aib71_ch3_x0y2, aib70_ch3_x0y2, aib69_ch3_x0y2,aib68_ch3_x0y2,
                                                   aib67_ch3_x0y2, aib66_ch3_x0y2, 1'b1,          aib64_ch3_x0y2,
                                                   aib63_ch3_x0y2, aib62_ch3_x0y2, 1'b1,          aib60_ch3_x0y2,
                                                   aib59_ch3_x0y2, aib58_ch3_x0y2, aib57_ch3_x0y2,aib56_ch3_x0y2,
                                                   aib55_ch3_x0y2, aib54_ch3_x0y2, aib53_ch3_x0y2,aib52_ch3_x0y2,
                                                   aib51_ch3_x0y2, aib50_ch3_x0y2, aib49_ch3_x0y2,aib48_ch3_x0y2,
                                                   aib47_ch3_x0y2, aib46_ch3_x0y2, aib45_ch3_x0y2,aib44_ch3_x0y2,
                                                   aib41_ch3_x0y2, aib40_ch3_x0y2, aib41_ch3_x0y2,aib40_ch3_x0y2,
                                                   aib19_ch3_x0y2, aib18_ch3_x0y2, aib17_ch3_x0y2,aib16_ch3_x0y2,
                                                   aib15_ch3_x0y2, aib14_ch3_x0y2, aib13_ch3_x0y2,aib12_ch3_x0y2,
                                                   aib11_ch3_x0y2, aib10_ch3_x0y2, aib9_ch3_x0y2, aib8_ch3_x0y2,
                                                   aib7_ch3_x0y2,  aib6_ch3_x0y2,  aib5_ch3_x0y2, aib4_ch3_x0y2,
                                                   aib3_ch3_x0y2,  aib2_ch3_x0y2,  aib1_ch3_x0y2, aib0_ch3_x0y2,
                                                   aib19_ch3_x0y2, aib18_ch3_x0y2, aib17_ch3_x0y2,aib16_ch3_x0y2,
                                                   aib15_ch3_x0y2, aib14_ch3_x0y2, aib13_ch3_x0y2,aib12_ch3_x0y2,
                                                   aib11_ch3_x0y2, aib10_ch3_x0y2, aib9_ch3_x0y2, aib8_ch3_x0y2,
                                                   aib7_ch3_x0y2,  aib6_ch3_x0y2,  aib5_ch3_x0y2, aib4_ch3_x0y2,
                                                   aib3_ch3_x0y2,  aib2_ch3_x0y2,  aib1_ch3_x0y2, aib0_ch3_x0y2}),
                    .io_aib_ch16                 ({aib95_ch4_x0y2, aib94_ch4_x0y2, 1'b1,         aib94_ch4_x0y2,
                                                   aib91_ch4_x0y2, aib90_ch4_x0y2, aib89_ch4_x0y2,aib88_ch4_x0y2,
                                                   aib87_ch4_x0y2, aib86_ch4_x0y2, aib85_ch4_x0y2,aib84_ch4_x0y2,
                                                   aib85_ch4_x0y2, aib84_ch4_x0y2, aib81_ch4_x0y2,aib80_ch4_x0y2,
                                                   aib79_ch4_x0y2, aib78_ch4_x0y2, aib77_ch4_x0y2,aib76_ch4_x0y2,
                                                   aib75_ch4_x0y2, aib74_ch4_x0y2, aib73_ch4_x0y2,aib72_ch4_x0y2,
                                                   aib71_ch4_x0y2, aib70_ch4_x0y2, aib69_ch4_x0y2,aib68_ch4_x0y2,
                                                   aib67_ch4_x0y2, aib66_ch4_x0y2, 1'b1,          aib64_ch4_x0y2,
                                                   aib63_ch4_x0y2, aib62_ch4_x0y2, 1'b1,          aib60_ch4_x0y2,
                                                   aib59_ch4_x0y2, aib58_ch4_x0y2, aib57_ch4_x0y2,aib56_ch4_x0y2,
                                                   aib55_ch4_x0y2, aib54_ch4_x0y2, aib53_ch4_x0y2,aib52_ch4_x0y2,
                                                   aib51_ch4_x0y2, aib50_ch4_x0y2, aib49_ch4_x0y2,aib48_ch4_x0y2,
                                                   aib47_ch4_x0y2, aib46_ch4_x0y2, aib45_ch4_x0y2,aib44_ch4_x0y2,
                                                   aib41_ch4_x0y2, aib40_ch4_x0y2, aib41_ch4_x0y2,aib40_ch4_x0y2,
                                                   aib19_ch4_x0y2, aib18_ch4_x0y2, aib17_ch4_x0y2,aib16_ch4_x0y2,
                                                   aib15_ch4_x0y2, aib14_ch4_x0y2, aib13_ch4_x0y2,aib12_ch4_x0y2,
                                                   aib11_ch4_x0y2, aib10_ch4_x0y2, aib9_ch4_x0y2, aib8_ch4_x0y2,
                                                   aib7_ch4_x0y2,  aib6_ch4_x0y2,  aib5_ch4_x0y2, aib4_ch4_x0y2,
                                                   aib3_ch4_x0y2,  aib2_ch4_x0y2,  aib1_ch4_x0y2, aib0_ch4_x0y2,
                                                   aib19_ch4_x0y2, aib18_ch4_x0y2, aib17_ch4_x0y2,aib16_ch4_x0y2,
                                                   aib15_ch4_x0y2, aib14_ch4_x0y2, aib13_ch4_x0y2,aib12_ch4_x0y2,
                                                   aib11_ch4_x0y2, aib10_ch4_x0y2, aib9_ch4_x0y2, aib8_ch4_x0y2,
                                                   aib7_ch4_x0y2,  aib6_ch4_x0y2,  aib5_ch4_x0y2, aib4_ch4_x0y2,
                                                   aib3_ch4_x0y2,  aib2_ch4_x0y2,  aib1_ch4_x0y2, aib0_ch4_x0y2}),
                    .io_aib_ch17                 ({aib95_ch5_x0y2, aib94_ch5_x0y2, 1'b1,         aib94_ch5_x0y2,
                                                   aib91_ch5_x0y2, aib90_ch5_x0y2, aib89_ch5_x0y2,aib88_ch5_x0y2,
                                                   aib87_ch5_x0y2, aib86_ch5_x0y2, aib85_ch5_x0y2,aib84_ch5_x0y2,
                                                   aib85_ch5_x0y2, aib84_ch5_x0y2, aib81_ch5_x0y2,aib80_ch5_x0y2,
                                                   aib79_ch5_x0y2, aib78_ch5_x0y2, aib77_ch5_x0y2,aib76_ch5_x0y2,
                                                   aib75_ch5_x0y2, aib74_ch5_x0y2, aib73_ch5_x0y2,aib72_ch5_x0y2,
                                                   aib71_ch5_x0y2, aib70_ch5_x0y2, aib69_ch5_x0y2,aib68_ch5_x0y2,
                                                   aib67_ch5_x0y2, aib66_ch5_x0y2, 1'b1,          aib64_ch5_x0y2,
                                                   aib63_ch5_x0y2, aib62_ch5_x0y2, 1'b1,          aib60_ch5_x0y2,
                                                   aib59_ch5_x0y2, aib58_ch5_x0y2, aib57_ch5_x0y2,aib56_ch5_x0y2,
                                                   aib55_ch5_x0y2, aib54_ch5_x0y2, aib53_ch5_x0y2,aib52_ch5_x0y2,
                                                   aib51_ch5_x0y2, aib50_ch5_x0y2, aib49_ch5_x0y2,aib48_ch5_x0y2,
                                                   aib47_ch5_x0y2, aib46_ch5_x0y2, aib45_ch5_x0y2,aib44_ch5_x0y2,
                                                   aib41_ch5_x0y2, aib40_ch5_x0y2, aib41_ch5_x0y2,aib40_ch5_x0y2,
                                                   aib19_ch5_x0y2, aib18_ch5_x0y2, aib17_ch5_x0y2,aib16_ch5_x0y2,
                                                   aib15_ch5_x0y2, aib14_ch5_x0y2, aib13_ch5_x0y2,aib12_ch5_x0y2,
                                                   aib11_ch5_x0y2, aib10_ch5_x0y2, aib9_ch5_x0y2, aib8_ch5_x0y2,
                                                   aib7_ch5_x0y2,  aib6_ch5_x0y2,  aib5_ch5_x0y2, aib4_ch5_x0y2,
                                                   aib3_ch5_x0y2,  aib2_ch5_x0y2,  aib1_ch5_x0y2, aib0_ch5_x0y2,
                                                   aib19_ch5_x0y2, aib18_ch5_x0y2, aib17_ch5_x0y2,aib16_ch5_x0y2,
                                                   aib15_ch5_x0y2, aib14_ch5_x0y2, aib13_ch5_x0y2,aib12_ch5_x0y2,
                                                   aib11_ch5_x0y2, aib10_ch5_x0y2, aib9_ch5_x0y2, aib8_ch5_x0y2,
                                                   aib7_ch5_x0y2,  aib6_ch5_x0y2,  aib5_ch5_x0y2, aib4_ch5_x0y2,
                                                   aib3_ch5_x0y2,  aib2_ch5_x0y2,  aib1_ch5_x0y2, aib0_ch5_x0y2}),
                    .io_aib_ch18                 ({aib95_ch0_x0y3, aib94_ch0_x0y3, 1'b1,         aib94_ch0_x0y3,
                                                   aib91_ch0_x0y3, aib90_ch0_x0y3, aib89_ch0_x0y3,aib88_ch0_x0y3,
                                                   aib87_ch0_x0y3, aib86_ch0_x0y3, aib85_ch0_x0y3,aib84_ch0_x0y3,
                                                   aib85_ch0_x0y3, aib84_ch0_x0y3, aib81_ch0_x0y3,aib80_ch0_x0y3,
                                                   aib79_ch0_x0y3, aib78_ch0_x0y3, aib77_ch0_x0y3,aib76_ch0_x0y3,
                                                   aib75_ch0_x0y3, aib74_ch0_x0y3, aib73_ch0_x0y3,aib72_ch0_x0y3,
                                                   aib71_ch0_x0y3, aib70_ch0_x0y3, aib69_ch0_x0y3,aib68_ch0_x0y3,
                                                   aib67_ch0_x0y3, aib66_ch0_x0y3, 1'b1,          aib64_ch0_x0y3,
                                                   aib63_ch0_x0y3, aib62_ch0_x0y3, 1'b1,          aib60_ch0_x0y3,
                                                   aib59_ch0_x0y3, aib58_ch0_x0y3, aib57_ch0_x0y3,aib56_ch0_x0y3,
                                                   aib55_ch0_x0y3, aib54_ch0_x0y3, aib53_ch0_x0y3,aib52_ch0_x0y3,
                                                   aib51_ch0_x0y3, aib50_ch0_x0y3, aib49_ch0_x0y3,aib48_ch0_x0y3,
                                                   aib47_ch0_x0y3, aib46_ch0_x0y3, aib45_ch0_x0y3,aib44_ch0_x0y3,
                                                   aib41_ch0_x0y3, aib40_ch0_x0y3, aib41_ch0_x0y3,aib40_ch0_x0y3,
                                                   aib19_ch0_x0y3, aib18_ch0_x0y3, aib17_ch0_x0y3,aib16_ch0_x0y3,
                                                   aib15_ch0_x0y3, aib14_ch0_x0y3, aib13_ch0_x0y3,aib12_ch0_x0y3,
                                                   aib11_ch0_x0y3, aib10_ch0_x0y3, aib9_ch0_x0y3, aib8_ch0_x0y3,
                                                   aib7_ch0_x0y3,  aib6_ch0_x0y3,  aib5_ch0_x0y3, aib4_ch0_x0y3,
                                                   aib3_ch0_x0y3,  aib2_ch0_x0y3,  aib1_ch0_x0y3, aib0_ch0_x0y3,
                                                   aib19_ch0_x0y3, aib18_ch0_x0y3, aib17_ch0_x0y3,aib16_ch0_x0y3,
                                                   aib15_ch0_x0y3, aib14_ch0_x0y3, aib13_ch0_x0y3,aib12_ch0_x0y3,
                                                   aib11_ch0_x0y3, aib10_ch0_x0y3, aib9_ch0_x0y3, aib8_ch0_x0y3,
                                                   aib7_ch0_x0y3,  aib6_ch0_x0y3,  aib5_ch0_x0y3, aib4_ch0_x0y3,
                                                   aib3_ch0_x0y3,  aib2_ch0_x0y3,  aib1_ch0_x0y3, aib0_ch0_x0y3}),
                    .io_aib_ch19                 ({aib95_ch1_x0y3, aib94_ch1_x0y3, 1'b1,         aib94_ch1_x0y3,
                                                   aib91_ch1_x0y3, aib90_ch1_x0y3, aib89_ch1_x0y3,aib88_ch1_x0y3,
                                                   aib87_ch1_x0y3, aib86_ch1_x0y3, aib85_ch1_x0y3,aib84_ch1_x0y3,
                                                   aib85_ch1_x0y3, aib84_ch1_x0y3, aib81_ch1_x0y3,aib80_ch1_x0y3,
                                                   aib79_ch1_x0y3, aib78_ch1_x0y3, aib77_ch1_x0y3,aib76_ch1_x0y3,
                                                   aib75_ch1_x0y3, aib74_ch1_x0y3, aib73_ch1_x0y3,aib72_ch1_x0y3,
                                                   aib71_ch1_x0y3, aib70_ch1_x0y3, aib69_ch1_x0y3,aib68_ch1_x0y3,
                                                   aib67_ch1_x0y3, aib66_ch1_x0y3, 1'b1,          aib64_ch1_x0y3,
                                                   aib63_ch1_x0y3, aib62_ch1_x0y3, 1'b1,          aib60_ch1_x0y3,
                                                   aib59_ch1_x0y3, aib58_ch1_x0y3, aib57_ch1_x0y3,aib56_ch1_x0y3,
                                                   aib55_ch1_x0y3, aib54_ch1_x0y3, aib53_ch1_x0y3,aib52_ch1_x0y3,
                                                   aib51_ch1_x0y3, aib50_ch1_x0y3, aib49_ch1_x0y3,aib48_ch1_x0y3,
                                                   aib47_ch1_x0y3, aib46_ch1_x0y3, aib45_ch1_x0y3,aib44_ch1_x0y3,
                                                   aib41_ch1_x0y3, aib40_ch1_x0y3, aib41_ch1_x0y3,aib40_ch1_x0y3,
                                                   aib19_ch1_x0y3, aib18_ch1_x0y3, aib17_ch1_x0y3,aib16_ch1_x0y3,
                                                   aib15_ch1_x0y3, aib14_ch1_x0y3, aib13_ch1_x0y3,aib12_ch1_x0y3,
                                                   aib11_ch1_x0y3, aib10_ch1_x0y3, aib9_ch1_x0y3, aib8_ch1_x0y3,
                                                   aib7_ch1_x0y3,  aib6_ch1_x0y3,  aib5_ch1_x0y3, aib4_ch1_x0y3,
                                                   aib3_ch1_x0y3,  aib2_ch1_x0y3,  aib1_ch1_x0y3, aib0_ch1_x0y3,
                                                   aib19_ch1_x0y3, aib18_ch1_x0y3, aib17_ch1_x0y3,aib16_ch1_x0y3,
                                                   aib15_ch1_x0y3, aib14_ch1_x0y3, aib13_ch1_x0y3,aib12_ch1_x0y3,
                                                   aib11_ch1_x0y3, aib10_ch1_x0y3, aib9_ch1_x0y3, aib8_ch1_x0y3,
                                                   aib7_ch1_x0y3,  aib6_ch1_x0y3,  aib5_ch1_x0y3, aib4_ch1_x0y3,
                                                   aib3_ch1_x0y3,  aib2_ch1_x0y3,  aib1_ch1_x0y3, aib0_ch1_x0y3}),
                    .io_aib_ch20                 ({aib95_ch2_x0y3, aib94_ch2_x0y3, 1'b1,         aib94_ch2_x0y3,
                                                   aib91_ch2_x0y3, aib90_ch2_x0y3, aib89_ch2_x0y3,aib88_ch2_x0y3,
                                                   aib87_ch2_x0y3, aib86_ch2_x0y3, aib85_ch2_x0y3,aib84_ch2_x0y3,
                                                   aib85_ch2_x0y3, aib84_ch2_x0y3, aib81_ch2_x0y3,aib80_ch2_x0y3,
                                                   aib79_ch2_x0y3, aib78_ch2_x0y3, aib77_ch2_x0y3,aib76_ch2_x0y3,
                                                   aib75_ch2_x0y3, aib74_ch2_x0y3, aib73_ch2_x0y3,aib72_ch2_x0y3,
                                                   aib71_ch2_x0y3, aib70_ch2_x0y3, aib69_ch2_x0y3,aib68_ch2_x0y3,
                                                   aib67_ch2_x0y3, aib66_ch2_x0y3, 1'b1,          aib64_ch2_x0y3,
                                                   aib63_ch2_x0y3, aib62_ch2_x0y3, 1'b1,          aib60_ch2_x0y3,
                                                   aib59_ch2_x0y3, aib58_ch2_x0y3, aib57_ch2_x0y3,aib56_ch2_x0y3,
                                                   aib55_ch2_x0y3, aib54_ch2_x0y3, aib53_ch2_x0y3,aib52_ch2_x0y3,
                                                   aib51_ch2_x0y3, aib50_ch2_x0y3, aib49_ch2_x0y3,aib48_ch2_x0y3,
                                                   aib47_ch2_x0y3, aib46_ch2_x0y3, aib45_ch2_x0y3,aib44_ch2_x0y3,
                                                   aib41_ch2_x0y3, aib40_ch2_x0y3, aib41_ch2_x0y3,aib40_ch2_x0y3,
                                                   aib19_ch2_x0y3, aib18_ch2_x0y3, aib17_ch2_x0y3,aib16_ch2_x0y3,
                                                   aib15_ch2_x0y3, aib14_ch2_x0y3, aib13_ch2_x0y3,aib12_ch2_x0y3,
                                                   aib11_ch2_x0y3, aib10_ch2_x0y3, aib9_ch2_x0y3, aib8_ch2_x0y3,
                                                   aib7_ch2_x0y3,  aib6_ch2_x0y3,  aib5_ch2_x0y3, aib4_ch2_x0y3,
                                                   aib3_ch2_x0y3,  aib2_ch2_x0y3,  aib1_ch2_x0y3, aib0_ch2_x0y3,
                                                   aib19_ch2_x0y3, aib18_ch2_x0y3, aib17_ch2_x0y3,aib16_ch2_x0y3,
                                                   aib15_ch2_x0y3, aib14_ch2_x0y3, aib13_ch2_x0y3,aib12_ch2_x0y3,
                                                   aib11_ch2_x0y3, aib10_ch2_x0y3, aib9_ch2_x0y3, aib8_ch2_x0y3,
                                                   aib7_ch2_x0y3,  aib6_ch2_x0y3,  aib5_ch2_x0y3, aib4_ch2_x0y3,
                                                   aib3_ch2_x0y3,  aib2_ch2_x0y3,  aib1_ch2_x0y3, aib0_ch2_x0y3}),
                    .io_aib_ch21                 ({aib95_ch3_x0y3, aib94_ch3_x0y3, 1'b1,         aib94_ch3_x0y3,
                                                   aib91_ch3_x0y3, aib90_ch3_x0y3, aib89_ch3_x0y3,aib88_ch3_x0y3,
                                                   aib87_ch3_x0y3, aib86_ch3_x0y3, aib85_ch3_x0y3,aib84_ch3_x0y3,
                                                   aib85_ch3_x0y3, aib84_ch3_x0y3, aib81_ch3_x0y3,aib80_ch3_x0y3,
                                                   aib79_ch3_x0y3, aib78_ch3_x0y3, aib77_ch3_x0y3,aib76_ch3_x0y3,
                                                   aib75_ch3_x0y3, aib74_ch3_x0y3, aib73_ch3_x0y3,aib72_ch3_x0y3,
                                                   aib71_ch3_x0y3, aib70_ch3_x0y3, aib69_ch3_x0y3,aib68_ch3_x0y3,
                                                   aib67_ch3_x0y3, aib66_ch3_x0y3, 1'b1,          aib64_ch3_x0y3,
                                                   aib63_ch3_x0y3, aib62_ch3_x0y3, 1'b1,          aib60_ch3_x0y3,
                                                   aib59_ch3_x0y3, aib58_ch3_x0y3, aib57_ch3_x0y3,aib56_ch3_x0y3,
                                                   aib55_ch3_x0y3, aib54_ch3_x0y3, aib53_ch3_x0y3,aib52_ch3_x0y3,
                                                   aib51_ch3_x0y3, aib50_ch3_x0y3, aib49_ch3_x0y3,aib48_ch3_x0y3,
                                                   aib47_ch3_x0y3, aib46_ch3_x0y3, aib45_ch3_x0y3,aib44_ch3_x0y3,
                                                   aib41_ch3_x0y3, aib40_ch3_x0y3, aib41_ch3_x0y3,aib40_ch3_x0y3,
                                                   aib19_ch3_x0y3, aib18_ch3_x0y3, aib17_ch3_x0y3,aib16_ch3_x0y3,
                                                   aib15_ch3_x0y3, aib14_ch3_x0y3, aib13_ch3_x0y3,aib12_ch3_x0y3,
                                                   aib11_ch3_x0y3, aib10_ch3_x0y3, aib9_ch3_x0y3, aib8_ch3_x0y3,
                                                   aib7_ch3_x0y3,  aib6_ch3_x0y3,  aib5_ch3_x0y3, aib4_ch3_x0y3,
                                                   aib3_ch3_x0y3,  aib2_ch3_x0y3,  aib1_ch3_x0y3, aib0_ch3_x0y3,
                                                   aib19_ch3_x0y3, aib18_ch3_x0y3, aib17_ch3_x0y3,aib16_ch3_x0y3,
                                                   aib15_ch3_x0y3, aib14_ch3_x0y3, aib13_ch3_x0y3,aib12_ch3_x0y3,
                                                   aib11_ch3_x0y3, aib10_ch3_x0y3, aib9_ch3_x0y3, aib8_ch3_x0y3,
                                                   aib7_ch3_x0y3,  aib6_ch3_x0y3,  aib5_ch3_x0y3, aib4_ch3_x0y3,
                                                   aib3_ch3_x0y3,  aib2_ch3_x0y3,  aib1_ch3_x0y3, aib0_ch3_x0y3}),
                    .io_aib_ch22                 ({aib95_ch4_x0y3, aib94_ch4_x0y3, 1'b1,         aib94_ch4_x0y3,
                                                   aib91_ch4_x0y3, aib90_ch4_x0y3, aib89_ch4_x0y3,aib88_ch4_x0y3,
                                                   aib87_ch4_x0y3, aib86_ch4_x0y3, aib85_ch4_x0y3,aib84_ch4_x0y3,
                                                   aib85_ch4_x0y3, aib84_ch4_x0y3, aib81_ch4_x0y3,aib80_ch4_x0y3,
                                                   aib79_ch4_x0y3, aib78_ch4_x0y3, aib77_ch4_x0y3,aib76_ch4_x0y3,
                                                   aib75_ch4_x0y3, aib74_ch4_x0y3, aib73_ch4_x0y3,aib72_ch4_x0y3,
                                                   aib71_ch4_x0y3, aib70_ch4_x0y3, aib69_ch4_x0y3,aib68_ch4_x0y3,
                                                   aib67_ch4_x0y3, aib66_ch4_x0y3, 1'b1,          aib64_ch4_x0y3,
                                                   aib63_ch4_x0y3, aib62_ch4_x0y3, 1'b1,          aib60_ch4_x0y3,
                                                   aib59_ch4_x0y3, aib58_ch4_x0y3, aib57_ch4_x0y3,aib56_ch4_x0y3,
                                                   aib55_ch4_x0y3, aib54_ch4_x0y3, aib53_ch4_x0y3,aib52_ch4_x0y3,
                                                   aib51_ch4_x0y3, aib50_ch4_x0y3, aib49_ch4_x0y3,aib48_ch4_x0y3,
                                                   aib47_ch4_x0y3, aib46_ch4_x0y3, aib45_ch4_x0y3,aib44_ch4_x0y3,
                                                   aib41_ch4_x0y3, aib40_ch4_x0y3, aib41_ch4_x0y3,aib40_ch4_x0y3,
                                                   aib19_ch4_x0y3, aib18_ch4_x0y3, aib17_ch4_x0y3,aib16_ch4_x0y3,
                                                   aib15_ch4_x0y3, aib14_ch4_x0y3, aib13_ch4_x0y3,aib12_ch4_x0y3,
                                                   aib11_ch4_x0y3, aib10_ch4_x0y3, aib9_ch4_x0y3, aib8_ch4_x0y3,
                                                   aib7_ch4_x0y3,  aib6_ch4_x0y3,  aib5_ch4_x0y3, aib4_ch4_x0y3,
                                                   aib3_ch4_x0y3,  aib2_ch4_x0y3,  aib1_ch4_x0y3, aib0_ch4_x0y3,
                                                   aib19_ch4_x0y3, aib18_ch4_x0y3, aib17_ch4_x0y3,aib16_ch4_x0y3,
                                                   aib15_ch4_x0y3, aib14_ch4_x0y3, aib13_ch4_x0y3,aib12_ch4_x0y3,
                                                   aib11_ch4_x0y3, aib10_ch4_x0y3, aib9_ch4_x0y3, aib8_ch4_x0y3,
                                                   aib7_ch4_x0y3,  aib6_ch4_x0y3,  aib5_ch4_x0y3, aib4_ch4_x0y3,
                                                   aib3_ch4_x0y3,  aib2_ch4_x0y3,  aib1_ch4_x0y3, aib0_ch4_x0y3}),
                    .io_aib_ch23                 ({aib95_ch5_x0y3, aib94_ch5_x0y3, 1'b1,         aib94_ch5_x0y3,
                                                   aib91_ch5_x0y3, aib90_ch5_x0y3, aib89_ch5_x0y3,aib88_ch5_x0y3,
                                                   aib87_ch5_x0y3, aib86_ch5_x0y3, aib85_ch5_x0y3,aib84_ch5_x0y3,
                                                   aib85_ch5_x0y3, aib84_ch5_x0y3, aib81_ch5_x0y3,aib80_ch5_x0y3,
                                                   aib79_ch5_x0y3, aib78_ch5_x0y3, aib77_ch5_x0y3,aib76_ch5_x0y3,
                                                   aib75_ch5_x0y3, aib74_ch5_x0y3, aib73_ch5_x0y3,aib72_ch5_x0y3,
                                                   aib71_ch5_x0y3, aib70_ch5_x0y3, aib69_ch5_x0y3,aib68_ch5_x0y3,
                                                   aib67_ch5_x0y3, aib66_ch5_x0y3, 1'b1,          aib64_ch5_x0y3,
                                                   aib63_ch5_x0y3, aib62_ch5_x0y3, 1'b1,          aib60_ch5_x0y3,
                                                   aib59_ch5_x0y3, aib58_ch5_x0y3, aib57_ch5_x0y3,aib56_ch5_x0y3,
                                                   aib55_ch5_x0y3, aib54_ch5_x0y3, aib53_ch5_x0y3,aib52_ch5_x0y3,
                                                   aib51_ch5_x0y3, aib50_ch5_x0y3, aib49_ch5_x0y3,aib48_ch5_x0y3,
                                                   aib47_ch5_x0y3, aib46_ch5_x0y3, aib45_ch5_x0y3,aib44_ch5_x0y3,
                                                   aib41_ch5_x0y3, aib40_ch5_x0y3, aib41_ch5_x0y3,aib40_ch5_x0y3,
                                                   aib19_ch5_x0y3, aib18_ch5_x0y3, aib17_ch5_x0y3,aib16_ch5_x0y3,
                                                   aib15_ch5_x0y3, aib14_ch5_x0y3, aib13_ch5_x0y3,aib12_ch5_x0y3,
                                                   aib11_ch5_x0y3, aib10_ch5_x0y3, aib9_ch5_x0y3, aib8_ch5_x0y3,
                                                   aib7_ch5_x0y3,  aib6_ch5_x0y3,  aib5_ch5_x0y3, aib4_ch5_x0y3,
                                                   aib3_ch5_x0y3,  aib2_ch5_x0y3,  aib1_ch5_x0y3, aib0_ch5_x0y3,
                                                   aib19_ch5_x0y3, aib18_ch5_x0y3, aib17_ch5_x0y3,aib16_ch5_x0y3,
                                                   aib15_ch5_x0y3, aib14_ch5_x0y3, aib13_ch5_x0y3,aib12_ch5_x0y3,
                                                   aib11_ch5_x0y3, aib10_ch5_x0y3, aib9_ch5_x0y3, aib8_ch5_x0y3,
                                                   aib7_ch5_x0y3,  aib6_ch5_x0y3,  aib5_ch5_x0y3, aib4_ch5_x0y3,
                                                   aib3_ch5_x0y3,  aib2_ch5_x0y3,  aib1_ch5_x0y3, aib0_ch5_x0y3}),
                    .io_aib_aux                  (AIB_AUX),
//                  .io_aib_aux                  (),
                    .io_aux_bg_ext_2k            (io_aux_bg_ext_2k),
	            .i_iocsr_rdy_aibaux          (top_io.i_adpt_hard_rst_n),
	            .i_aibaux_por_vccl_ovrd      (1'b1),      
                    .i_aibaux_ctrl_bus0          (32'b0), 
//                  .i_aibaux_ctrl_bus1          (32'h805001e0),  //observe oosc dft[12:0] 
                    .i_aibaux_ctrl_bus1          (32'h00500020),  //observe oosc dft[12:0] 
                    .i_aibaux_ctrl_bus2          (32'b0), 
                    .i_aibaux_osc_fuse_trim      (10'b0), 
//                  .i_osc_bypclk                (i_osc_clk),  
                    .i_osc_bypclk                (1'b0),  
                    .o_aibaux_osc_clk            (),      
                    .i_scan_clk                  (1'b0), 
                    .i_test_clk_125m             (1'b0), 
                    .i_test_clk_1g               (1'b0), 
                    .i_test_clk_250m             (1'b0), 
                    .i_test_clk_500m             (1'b0), 
                    .i_test_clk_62m              (1'b0), 	      
                    .i_test_c3adapt_scan_in      ({24*17{1'b0}}),
//                  .i_test_c3adapt_tcb_static_common (60'h010_8421_0842_1000),
                    .i_test_c3adapt_tcb_static_common (60'h050_8421_0842_1000),
	            .o_test_c3adapt_scan_out     (),
                    .i_jtag_clkdr                (1'b0),   
                    .i_jtag_clksel               (1'b0),   
                    .i_jtag_intest               (1'b0),   
                    .i_jtag_mode                 (1'b0),   
                    .i_jtag_rstb_en              (1'b0),   
                    .i_jtag_rstb                 (1'b0),   
                    .i_jtag_weakpdn              (1'b0),   
                    .i_jtag_weakpu               (1'b0), 	      
                    .i_jtag_tx_scan              (1'b0),
                    .i_jtag_tx_scanen            (1'b0),
                    .i_aibdft2osc                ({1'b0, 1'b1, i_rx_pma_div2_clk}),
                    .o_aibdft2osc                (),
                    .o_last_bs_out               (),
                    .o_por                       (),
                    .o_osc_monitor               (),
                    .i_aux_atpg_mode_n           (1'b1),  //FIXME
                    .i_aux_atpg_pipeline_global_en (1'b0),  //FIXME
                    .i_aux_atpg_rst_n            (1'b1),  //FIXME
                    .i_aux_atpg_scan_clk         (1'b0),
                    .i_aux_atpg_scan_in          (1'b0),
                    .i_aux_atpg_scan_shift_n     (1'b1),  //FIXME
                    .o_aux_atpg_scan_out         ()    	      
               );

    
endmodule 

