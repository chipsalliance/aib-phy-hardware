// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. 
// Library - aibnd_lib, Cell - aibnd_txdatapath_tx, View - schematic
// LAST TIME SAVED: Jul  7 15:46:47 2015
// NETLIST TIME: Jul  8 13:09:52 2015
// `timescale 1ns / 1ns 

module aibnd_txdatapath_tx ( async_dat_outpdir1_1, dcc_done,
     dft_rx_clk, iasyncdata_oshared2, idat0_outpdir6, idat0_poutp18,
     idat1_poutp18, idataselb_oshared2, idataselb_outpdir1_1,
     idataselb_outpdir6, idataselb_poutp18, iddren_poutp18,
     ilaunch_clk_poutp18, irxen_chain2, irxen_inpclk3, irxen_inpdir3,
     irxen_inpshared0, irxen_inpshared4, irxen_ptxclkin,
     itxen_oshared2, itxen_outpdir1_1, itxen_outpdir6, itxen_poutp18,
     jtag_clkdr_inpclk0n, jtag_clkdr_inpshared0, jtag_clkdr_inpshared4,
     jtag_clkdr_oshared2, jtag_clkdr_out_chain2,
     jtag_clkdr_out_inpclk3, jtag_clkdr_out_inpdir3,
     jtag_clkdr_out_outpdir1_1, jtag_clkdr_out_outpdir6,
     jtag_clkdr_out_poutp18, jtag_clkdr_ptxclkin, jtag_clkdr_ptxclkinn,
     jtag_rx_scan_inpclk0n, jtag_rx_scan_inpshared0,
     jtag_rx_scan_inpshared4, jtag_rx_scan_oshared2,
     jtag_rx_scan_out_inpclk3, jtag_rx_scan_out_inpdir3,
     jtag_rx_scan_out_outpdir1_1, jtag_rx_scan_out_outpdir6,
     jtag_rx_scan_out_poutp18, jtag_rx_scan_ptxclkin,
     jtag_rx_scan_ptxclkinn, jtag_scan_out_chain2, oaibdftcore2dll,
     oaibdftdll2core, oclk_inpclk3, oclkb_inpclk3, oclkn_inpclk3,
     oclkn_outpdir4_1, odat0_inpdir0, odat1_inpdir0, odat_async,
     odat_async_oshared1, odat_async_pout0, odirectin_data,
     odirectin_data_out0_chain2, out_rx_fast_clk, scan_out,
     shift_en_inpclk0n, shift_en_inpclk3, shift_en_inpdir3,
     shift_en_inpshared0, shift_en_inpshared4, shift_en_oshared2,
     shift_en_out_chain2, shift_en_outpdir1_1, shift_en_outpdir6,
     shift_en_poutp18, shift_en_ptxclkin, shift_en_ptxclkinn,
     iopad_async_in, iopad_async_out, iopad_clkn, iopad_clkp,
     iopad_dat, iopad_direct_input, iopad_directinclkn,
     iopad_directinclkp, iopad_directout, async_dat_outpclk1_1,
     async_dat_outpdir0_1, avmm_sync_rstb, clkdr_xr1l, clkdr_xr1r,
     clkdr_xr2l, clkdr_xr2r, clkdr_xr3l, clkdr_xr3r, clkdr_xr4l,
     clkdr_xr4r, clkdr_xr5l, clkdr_xr5r, clkdr_xr6l, clkdr_xr6r,
     clkdr_xr7l, clkdr_xr7r, clkdr_xr8l, clkdr_xr8r, csr_reg,
     dcc_dft_nrst, dcc_dft_nrst_coding, dcc_dft_up, dcc_req,
     dll_csr_reg6, iaibdftcore2dll, iasyncdata, iclkin_dist_pinp0,
     idat0, idat0_clkn, idat0_clkp, idat0_in0_dout_clkp, idat0_voutp00,
     idat0_voutp01, idat1, idat1_clkn, idat1_clkp, idat1_in0_dout_clkp,
     idat1_voutp00, idat1_voutp01, idata0_ssrdout, idata0_ssrldout,
     idata1_ssrdout, idata1_ssrldout, idataselb,
     idataselb_in0_dout_clkp, idataselb_outpclk1_1,
     idataselb_outpdir0_1, idataselb_ssrdout, idataselb_ssrldout,
     idataselb_voutp00, idataselb_voutp01, iddren, idirectout_data,
     idll_dll2core, idll_entest, ilaunch_clk_in0_dout_clkp,
     ilaunch_clk_ssrdout, ilaunch_clk_ssrldout, ilaunch_clk_voutp00,
     ilaunch_clk_voutp01, indrv_r12, indrv_r34, indrv_r56, ipdrv_r12,
     ipdrv_r34, ipdrv_r56, irxen_in_chain2, irxen_inpclk6,
     irxen_inpdir2, irxen_pinp0, irxen_r0, irxen_r1, irxen_r2,
     istrbclk_pinp0, itxen, itxen_in0_dout_clkp, itxen_outpclk1_1,
     itxen_outpdir0_1, itxen_ssrdout, itxen_ssrldout, itxen_voutp00,
     itxen_voutp01, jtag_clkdr_in_chain2, jtag_clkdr_in_ssrdout,
     jtag_clkdr_in_ssrldout, jtag_clkdr_inpclk1n, jtag_clkdr_inpclk6,
     jtag_clkdr_out_diin_clkp, jtag_clkdr_out_directin2,
     jtag_clkdr_outpclk1_1, jtag_clkdr_outpdir0_1, jtag_clkdr_pinp0,
     jtag_clkdr_voutp00, jtag_clkdr_voutp01, jtag_clksel, jtag_intest,
     jtag_mode_in, jtag_rstb, jtag_rstb_en, jtag_rx_scan_in_ssrdout,
     jtag_rx_scan_in_ssrldout, jtag_rx_scan_inpclk1n,
     jtag_rx_scan_inpclk6, jtag_rx_scan_out_diin_clkp,
     jtag_rx_scan_out_directin2, jtag_rx_scan_outpclk1_1,
     jtag_rx_scan_outpdir0_1, jtag_rx_scan_voutp00,
     jtag_rx_scan_voutp01, jtag_scan_in_chain2, jtag_scan_pinp0,
     jtag_tx_scanen_in, jtag_weakpdn, jtag_weakpu, oclk_inpdir2,
     oclk_srclkout, oclkb_inpdir2, oclkb_srclkout, oclkn_inpdir4,
     odat_async_chain2, odat_async_fsrdin, odat_async_inpclk1,
     odat_async_inpclk4, output_buffer_clk, output_rstb,
     pipeline_global_en, poutp_dig_rstb, rb_clkdiv, rb_dcc_byp,
     rb_dcc_byp_dprio, // Mod : Added new port 
     rb_dcc_dft, rb_dcc_dft_sel, rb_dcc_dll_dft_sel, rb_dcc_en,
     rb_dcc_en_dprio, //Mod : Added new port
     rb_dcc_manual_dn, rb_dcc_manual_mode, 
     rb_dcc_manual_mode_dprio, // Mod : Added new port  
     rb_dcc_manual_up,
     rb_dcc_test_clk_pll_en_n, rb_half_code, rb_selflock,
     rshift_en_dirclkn, rshift_en_dirclkp, rshift_en_drx,
     rshift_en_dtx, rshift_en_poutp, rshift_en_rx, rshift_en_tx,
     rshift_en_txferclkout, rshift_en_txferclkoutn, scan_clk_in,
     scan_in, scan_mode_n, scan_rst_n, scan_shift_n,
     shift_en_in_chain2, shift_en_inpclk1n, shift_en_inpclk6,
     shift_en_inpdir2, shift_en_outpclk0, shift_en_outpclk1_1,
     shift_en_outpdir0_1, shift_en_pinp0, shift_en_ssrdout,
     shift_en_ssrldout, shift_en_voutp00, shift_en_voutp01, vccl_aibnd,
     vssl_aibnd );

output  async_dat_outpdir1_1, dcc_done, dft_rx_clk,
     iasyncdata_oshared2, idat0_outpdir6, idat0_poutp18, idat1_poutp18,
     idataselb_oshared2, idataselb_outpdir1_1, idataselb_outpdir6,
     idataselb_poutp18, iddren_poutp18, ilaunch_clk_poutp18,
     itxen_oshared2, itxen_outpdir1_1, itxen_outpdir6, itxen_poutp18,
     jtag_clkdr_inpclk0n, jtag_clkdr_inpshared0, jtag_clkdr_inpshared4,
     jtag_clkdr_oshared2, jtag_clkdr_out_chain2,
     jtag_clkdr_out_inpclk3, jtag_clkdr_out_inpdir3,
     jtag_clkdr_out_outpdir1_1, jtag_clkdr_out_outpdir6,
     jtag_clkdr_out_poutp18, jtag_clkdr_ptxclkin, jtag_clkdr_ptxclkinn,
     jtag_rx_scan_inpclk0n, jtag_rx_scan_inpshared0,
     jtag_rx_scan_inpshared4, jtag_rx_scan_oshared2,
     jtag_rx_scan_out_inpclk3, jtag_rx_scan_out_inpdir3,
     jtag_rx_scan_out_outpdir1_1, jtag_rx_scan_out_outpdir6,
     jtag_rx_scan_out_poutp18, jtag_rx_scan_ptxclkin,
     jtag_rx_scan_ptxclkinn, jtag_scan_out_chain2, oclk_inpclk3,
     oclkb_inpclk3, oclkn_inpclk3, oclkn_outpdir4_1, odat0_inpdir0,
     odat1_inpdir0, odat_async_oshared1, odat_async_pout0,
     odirectin_data_out0_chain2, scan_out, shift_en_inpclk0n,
     shift_en_inpclk3, shift_en_inpdir3, shift_en_inpshared0,
     shift_en_inpshared4, shift_en_oshared2, shift_en_out_chain2,
     shift_en_outpdir1_1, shift_en_outpdir6, shift_en_poutp18,
     shift_en_ptxclkin, shift_en_ptxclkinn;

inout  iopad_clkn, iopad_clkp;

input  async_dat_outpclk1_1, async_dat_outpdir0_1, avmm_sync_rstb,
     clkdr_xr1l, clkdr_xr1r, clkdr_xr2l, clkdr_xr2r, clkdr_xr3l,
     clkdr_xr3r, clkdr_xr4l, clkdr_xr4r, clkdr_xr5l, clkdr_xr5r,
     clkdr_xr6l, clkdr_xr6r, clkdr_xr7l, clkdr_xr7r, clkdr_xr8l,
     clkdr_xr8r, dcc_dft_nrst, dcc_dft_nrst_coding, dcc_dft_up,
     dcc_req, dll_csr_reg6, iclkin_dist_pinp0, idat0_clkn, idat0_clkp,
     idat0_in0_dout_clkp, idat0_voutp00, idat0_voutp01, idat1_clkn,
     idat1_clkp, idat1_in0_dout_clkp, idat1_voutp00, idat1_voutp01,
     idata0_ssrdout, idata0_ssrldout, idata1_ssrdout, idata1_ssrldout,
     idataselb_in0_dout_clkp, idataselb_outpclk1_1,
     idataselb_outpdir0_1, idataselb_ssrdout, idataselb_ssrldout,
     idataselb_voutp00, idataselb_voutp01, iddren, idll_entest,
     ilaunch_clk_in0_dout_clkp, ilaunch_clk_ssrdout,
     ilaunch_clk_ssrldout, ilaunch_clk_voutp00, ilaunch_clk_voutp01,
     istrbclk_pinp0, itxen_in0_dout_clkp, itxen_outpclk1_1,
     itxen_outpdir0_1, itxen_ssrdout, itxen_ssrldout, itxen_voutp00,
     itxen_voutp01, jtag_clkdr_in_chain2, jtag_clkdr_in_ssrdout,
     jtag_clkdr_in_ssrldout, jtag_clkdr_inpclk1n, jtag_clkdr_inpclk6,
     jtag_clkdr_out_diin_clkp, jtag_clkdr_out_directin2,
     jtag_clkdr_outpclk1_1, jtag_clkdr_outpdir0_1, jtag_clkdr_pinp0,
     jtag_clkdr_voutp00, jtag_clkdr_voutp01, jtag_clksel, jtag_intest,
     jtag_mode_in, jtag_rstb, jtag_rstb_en, jtag_rx_scan_in_ssrdout,
     jtag_rx_scan_in_ssrldout, jtag_rx_scan_inpclk1n,
     jtag_rx_scan_inpclk6, jtag_rx_scan_out_diin_clkp,
     jtag_rx_scan_out_directin2, jtag_rx_scan_outpclk1_1,
     jtag_rx_scan_outpdir0_1, jtag_rx_scan_voutp00,
     jtag_rx_scan_voutp01, jtag_scan_in_chain2, jtag_scan_pinp0,
     jtag_tx_scanen_in, jtag_weakpdn, jtag_weakpu, oclk_inpdir2,
     oclk_srclkout, oclkb_inpdir2, oclkb_srclkout, oclkn_inpdir4,
     odat_async_chain2, odat_async_fsrdin, odat_async_inpclk1,
     odat_async_inpclk4, output_buffer_clk, output_rstb,
     pipeline_global_en, poutp_dig_rstb, rb_dcc_byp, 
     rb_dcc_byp_dprio, // Mod : Added new port 
     rb_dcc_dft,
     rb_dcc_dft_sel, rb_dcc_dll_dft_sel, rb_dcc_en, 
     rb_dcc_en_dprio, // Mod : Added new port
     rb_dcc_manual_mode,
     rb_dcc_manual_mode_dprio, // Mod : Added new port 
     rb_dcc_test_clk_pll_en_n, rb_half_code, rb_selflock,
     rshift_en_txferclkout, rshift_en_txferclkoutn, scan_clk_in,
     scan_in, scan_mode_n, scan_rst_n, scan_shift_n,
     shift_en_in_chain2, shift_en_inpclk1n, shift_en_inpclk6,
     shift_en_inpdir2, shift_en_outpclk0, shift_en_outpclk1_1,
     shift_en_outpdir0_1, shift_en_pinp0, shift_en_ssrdout,
     shift_en_ssrldout, shift_en_voutp00, shift_en_voutp01, vccl_aibnd,
     vssl_aibnd;

output [2:0]  irxen_chain2;
output [2:0]  irxen_inpclk3;
output [12:0]  oaibdftdll2core;
output [2:0]  irxen_inpdir3;
output [2:0]  irxen_inpshared0;
output [2:0]  irxen_ptxclkin;
output [2:0]  oaibdftcore2dll;
output [2:0]  odirectin_data;
output [2:0]  irxen_inpshared4;
output [4:0]  odat_async;
output [1:0]  out_rx_fast_clk;

inout [2:0]  iopad_direct_input;
inout [1:0]  iopad_directinclkp;
inout [1:0]  iopad_directinclkn;
inout [2:0]  iopad_async_out;
inout [4:0]  iopad_async_in;
inout [3:0]  iopad_directout;
inout [19:0]  iopad_dat;

input [1:0]  indrv_r34;
input [1:0]  ipdrv_r34;
input [2:0]  irxen_inpdir2;
input [12:0]  idll_dll2core;
input [1:0]  ipdrv_r12;
input [2:0]  irxen_r0;
input [1:0]  indrv_r12;
input [1:0]  ipdrv_r56;
input [1:0]  indrv_r56;
input [2:0]  irxen_pinp0;
input [2:0]  irxen_in_chain2;
input [1:0]  rshift_en_dirclkn;
input [2:0]  irxen_inpclk6;
input [2:0]  iaibdftcore2dll;
input [1:0]  rshift_en_dirclkp;
input [51:0]  csr_reg;
input [2:0]  irxen_r1;
input [2:0]  rshift_en_drx;
input [4:0]  rb_dcc_manual_up;
input [4:0]  rb_dcc_manual_dn;
input [2:0]  iasyncdata;
input [2:0]  irxen_r2;
input [3:0]  rshift_en_rx;
input [2:0]  rb_clkdiv;
input [3:0]  rshift_en_tx;
input [3:0]  rshift_en_dtx;
input [3:0]  idirectout_data;
input [19:0]  rshift_en_poutp;
input [3:0]  idataselb;
input [3:0]  itxen;
input [19:0]  idat1;
input [19:0]  idat0;

wire output_buffer_clk, outbuf_clk_buf, rb_dcc_dll_dft_sel, dcc_scan_out, scan_out, clk_mimic0, clk_mimic0_buf, clk_mimic1, clk_mimic1_buf, gated_clk_mimic1, dft_rx_clk, dll_csr_reg6, nc_clk_repb, clk_rep, nc_clk_mimic, clk_mimic; // Conversion Sript Generated

wire out_rx_fast_clk0_buf;
wire nc_out_rx_fast_clk0_io;

// Buses in the design

wire  [1:1]  ncdtx_oclkb_aib;

wire  [0:0]  drx_oclk_aib;

wire  [0:12]  mux_dft_dll2core;

wire  [0:12]  buf_dcc2core;

wire  [2:0]  oaibdftcore2dcc;

wire  [4:4]  ncrx_oclk;

wire  [0:0]  ncdrx_odat0_aib;

wire  [0:1]  ncout_rx_fast_clkn;

wire  [0:1]  ncout_rx_fast_clknb;

wire  [0:1]  nc_rxodat0_clkn;

wire  [0:1]  nc_rxodat1_clkn;

wire  [0:1]  nc_rxodat_async_clkn;

wire  [0:1]  nc_rxpd_data_clkn;

wire  [0:1]  out_rx_fast_clkb;

wire  [0:1]  nc_rxodat0_clkp;

wire  [0:1]  nc_rxodat1_clkp;

wire  [0:1]  nc_rxodat_async_clkp;

wire  [0:1]  nc_rxpd_data_clkp;

wire  [1:1]  ncdrx_oclk_aib;

wire  [1:1]  ncdrx_oclkb_aib;

wire  [0:2]  ncdrx_oclk;

wire  [0:2]  ncdrx_oclkb;

wire  [0:2]  ncdrx_odat0;

wire  [0:2]  ncdrx_odat1;

wire  [0:2]  ncdrx_pd_data;

wire  [2:2]  ncdrx_odat1_aib;

wire  [0:2]  nctx_odat_async;

wire  [0:12]  buf_dll2core;

wire  [0:0]  drx_oclkb_aib;

wire  [4:4]  ncrx_oclk_aib;

wire  [4:4]  ncrx_oclkb_aib;

wire  [0:2]  ncdrx_odat_async_aib;

wire  [0:2]  nctx_oclkn;

wire  [0:2]  nctx_oclk;

wire  [0:2]  nctx_oclkb;

wire  [0:2]  nctx_odat0;

wire  [0:2]  nctx_odat1;

wire  [0:2]  nctx_pd_data;

wire  [0:2]  nctx_oclk_aib;

wire  [0:2]  nctx_oclkb_aib;

wire  [0:2]  nctx_odat0_aib;

wire  [0:2]  nctx_odat1_aib;

wire  [0:2]  nctx_pd_data_aib;

wire  [0:11]  tx_launch_clk_l;

wire  [0:4]  ncrx_odat0_aib;

wire  [0:4]  ncrx_odat1_aib;

wire  [0:4]  ncrx_pd_data_aib;

wire  [0:4]  ncrx_oclkb;

wire  [0:4]  ncrx_odat0;

wire  [0:4]  ncrx_odat1;

wire  [0:4]  ncrx_pd_data;

wire  [3:3]  ncdtx_oclk_aib;

wire  [0:3]  ncrx_odat_async_aib;

wire  [2:3]  ncdtx_oclkn;

wire  [0:2]  ncdrx_pd_data_aib;

wire  [0:11]  tx_launch_clk_r;

wire  [0:3]  ncdtx_oclk;

wire  [0:3]  ncdtx_oclkb;

wire  [0:3]  ncdtx_odat0;

wire  [0:3]  ncdtx_odat1;

wire  [0:3]  ncdtx_odat_async;

wire  [0:3]  ncdtx_pd_data;

wire  [0:3]  ncdtx_odat0_aib;

wire  [0:3]  ncdtx_odat1_aib;

wire  [0:1]  ncdtx_odat_async_aib;

wire  [0:3]  ncdtx_pd_data_aib;

wire  [12:0]  odcc_dll2core;

wire  [0:19]  nc_oclkn_pout;

wire  [0:19]  nc_oclkb_aib_pout;

wire  [0:19]  nc_odat1_aib_pout;

wire  [0:19]  nc_pd_data_aib_pout;

wire  [0:19]  nc_oclk;

wire  [0:19]  nc_oclkb;

wire  [0:19]  nc_odat1;

wire  [0:19]  nc_odat0_aib_pout;

wire  [1:19]  nc_odat_async_aib_pout;

wire  [0:19]  nc_odat_async;

wire  [0:19]  nc_odat0;

wire  [0:19]  nc_oclk_aib_pout;

wire  [0:19]  nc_pd_data;


// specify 
//     specparam CDS_LIBNAME  = "aibnd_lib";
//     specparam CDS_CELLNAME = "aibnd_txdatapath_tx";
//     specparam CDS_VIEWNAME = "schematic";
// endspecify

aibnd_clktree  xclktree ( //.vcc_aibnd(vccl_aibnd),
     //.vss_aibnd(vssl_aibnd), 
	 .lstrbclk_r_11(tx_launch_clk_r[11]),
     .lstrbclk_r_10(tx_launch_clk_r[10]),
     .lstrbclk_l_11(tx_launch_clk_l[11]), .lstrbclk_mimic2(clk_mimic),
     .lstrbclk_mimic1(clk_mimic1), .lstrbclk_mimic0(clk_mimic0),
     .lstrbclk_l_10(tx_launch_clk_l[10]),
     .lstrbclk_r_9(tx_launch_clk_r[9]),
     .lstrbclk_r_8(tx_launch_clk_r[8]),
     .lstrbclk_r_7(tx_launch_clk_r[7]),
     .lstrbclk_r_6(tx_launch_clk_r[6]),
     .lstrbclk_r_5(tx_launch_clk_r[5]),
     .lstrbclk_r_4(tx_launch_clk_r[4]),
     .lstrbclk_r_3(tx_launch_clk_r[3]),
     .lstrbclk_r_2(tx_launch_clk_r[2]),
     .lstrbclk_r_1(tx_launch_clk_r[1]),
     .lstrbclk_r_0(tx_launch_clk_r[0]),
     .lstrbclk_l_0(tx_launch_clk_l[0]),
     .lstrbclk_l_1(tx_launch_clk_l[1]),
     .lstrbclk_l_2(tx_launch_clk_l[2]),
     .lstrbclk_l_3(tx_launch_clk_l[3]),
     .lstrbclk_l_4(tx_launch_clk_l[4]),
     .lstrbclk_l_5(tx_launch_clk_l[5]),
     .lstrbclk_l_6(tx_launch_clk_l[6]),
     .lstrbclk_l_7(tx_launch_clk_l[7]),
     .lstrbclk_l_8(tx_launch_clk_l[8]),
     .lstrbclk_l_9(tx_launch_clk_l[9]), .lstrbclk_rep(clk_rep),
     .clkin(clktree_in));
aibnd_buffx1_top xasyncrx3 ( .idata1_in1_jtag_out(nc_idat1_async_in3),
     .async_dat_in1_jtag_out(nc_async_dat_async_in3),
     .idata0_in1_jtag_out(nc_idat0_async_in3),
     .jtag_clkdr_outn(jtag_clkdr_outn_inpshared3),
     .prev_io_shift_en(shift_en_ssrldout), .anlg_rstb(output_rstb),
     .pd_data_aib(ncrx_pd_data_aib[3]), .oclk_out(odat_async[3]),
     .oclkb_out(ncrx_oclkb[3]), .odat0_out(ncrx_odat0[3]),
     .odat1_out(ncrx_odat1[3]), .odat_async_out(ncrx_async_data_out3),
     .pd_data_out(ncrx_pd_data[3]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(vssl_aibnd),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(idata0_ssrldout), .idata1_in0(vssl_aibnd),
     .idata1_in1(idata1_ssrldout), .idataselb_in0(vssl_aibnd),
     .idataselb_in1(idataselb_ssrldout), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(ilaunch_clk_ssrldout),
     .ilpbk_dat_in0(vssl_aibnd), .ilpbk_dat_in1(vssl_aibnd),
     .ilpbk_en_in0(vssl_aibnd), .ilpbk_en_in1(vssl_aibnd),
     .indrv_in0({vssl_aibnd, vssl_aibnd}), .indrv_in1(indrv_r34[1:0]),
     .ipdrv_in0({vssl_aibnd, vssl_aibnd}), .ipdrv_in1(ipdrv_r34[1:0]),
     .irxen_in0({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(vssl_aibnd), .itxen_in1(itxen_ssrldout),
     .oclk_in1(vssl_aibnd), .odat_async_aib(ncrx_odat_async_aib[3]),
     .oclkb_in1(vssl_aibnd), .jtag_clksel(jtag_clksel),
     .odat0_in1(vssl_aibnd), .vssl_aibnd(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_tx[3]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(avmm_sync_rstb), .jtag_clkdr_out(jtag_clkdr_async_in3),
     .jtag_intest(jtag_intest), .odat1_aib(ncrx_odat1_aib[3]),
     .jtag_rx_scan_out(jtag_rx_scan_async_in3),
     .odat0_aib(ncrx_odat0_aib[3]), .oclk_aib(ncrx_oclk_aib3),
     .last_bs_out(nc_last_bs_out_diro3), .vccl_aibnd(vccl_aibnd),
     .oclkb_aib(ncrx_oclkb_aib3), .jtag_clkdr_in(clkdr_xr4r),
     .jtag_rstb_en(jtag_rstb_en), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_in_ssrldout),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_async_in[3]), .oclkn(oclkn_inpshared3),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xasyncrx1 ( .idata1_in1_jtag_out(nc_idat1_async_in1),
     .async_dat_in1_jtag_out(nc_async_dat_async_in1),
     .idata0_in1_jtag_out(nc_idat0_async_in1),
     .jtag_clkdr_outn(jtag_clkdr_outn_inpshared1),
     .prev_io_shift_en(rshift_en_tx[3]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(output_rstb), .pd_data_aib(ncrx_pd_data_aib[1]),
     .oclk_out(odat_async[1]), .oclkb_out(ncrx_oclkb[1]),
     .odat0_out(ncrx_odat0[1]), .odat1_out(ncrx_odat1[1]),
     .odat_async_out(ncrx_async_data_out1),
     .pd_data_out(ncrx_pd_data[1]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(vssl_aibnd),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vssl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(ncrx_odat_async_aib[1]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_tx[1]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(output_rstb), .jtag_clkdr_out(jtag_clkdr_async_in1),
     .odat1_aib(ncrx_odat1_aib[1]),
     .jtag_rx_scan_out(jtag_rx_scan_async_in1),
     .odat0_aib(ncrx_odat0_aib[1]), .oclk_aib(ncrx_oclk_aib1),
     .last_bs_out(nc_last_bs_out_diro1), .oclkb_aib(ncrx_oclkb_aib1),
     .jtag_clkdr_in(clkdr_xr4r), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_async_in3),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_async_in[1]), .oclkn(oclkn_inpshared1),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top x455 ( .idata1_in1_jtag_out(idat1_poutp9),
     .async_dat_in1_jtag_out(nc_async_dat_poutp9),
     .idata0_in1_jtag_out(idat0_poutp9),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp9),
     .prev_io_shift_en(rshift_en_poutp[7]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_pout[9]), .oclk_out(nc_oclk[9]),
     .oclkb_out(nc_oclkb[9]), .odat0_out(nc_odat0[9]),
     .odat1_out(nc_odat1[9]), .odat_async_out(nc_odat_async[9]),
     .pd_data_out(nc_pd_data[9]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp9),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[9]),
     .idata0_in1(idat0_poutp7), .idata1_in0(idat1[9]),
     .idata1_in1(idat1_poutp7), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[0]), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk_r[4]),
     .ilaunch_clk_in1(tx_launch_clk_r[4]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp9), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[9]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[9]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_poutp9),
     .odat1_aib(nc_odat1_aib_pout[9]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp9),
     .odat0_aib(nc_odat0_aib_pout[9]), .oclk_aib(nc_oclk_aib_pout[9]),
     .last_bs_out(nc_last_bs_out_poutp9),
     .oclkb_aib(nc_oclkb_aib_pout[9]), .jtag_clkdr_in(clkdr_xr6r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp7),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[9]), .oclkn(nc_oclkn_pout[9]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top x454 ( .idata1_in1_jtag_out(idata1_in1_clkn),
     .async_dat_in1_jtag_out(nc_async_dat_clkn),
     .idata0_in1_jtag_out(idata0_in1_clkn),
     .jtag_clkdr_outn(jtag_clkdr_outn_clkn),
     .prev_io_shift_en(rshift_en_poutp[9]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_txferclkoutn),
     .oclk_out(nc_oclk_clkn), .oclkb_out(nc_oclkb_clkn),
     .odat0_out(nc_odat0_clkn), .odat1_out(nc_odat1_clkn),
     .odat_async_out(nc_odat_async_clkn),
     .pd_data_out(nc_pd_data_clkn), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_clkn),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0_clkn),
     .idata0_in1(idat0_poutp9), .idata1_in0(idat1_clkn),
     .idata1_in1(idat1_poutp9), .idataselb_in0(idataselb[1]),
     .idataselb_in1(idataselb[0]), .iddren_in0(vccl_aibnd),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk_r[8]),
     .ilaunch_clk_in1(tx_launch_clk_r[8]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_clkn), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[1]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_txferclkoutn),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_txferclkoutn), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_clkn),
     .odat1_aib(nc_odat1_aib_txferclkoutn),
     .jtag_rx_scan_out(jtag_rx_scan_out_clkn),
     .odat0_aib(nc_odat0_aib_txferclkoutn),
     .oclk_aib(nc_oclk_aib_txferclkoutn),
     .last_bs_out(nc_last_bs_out_txferclkoutn),
     .oclkb_aib(nc_oclkb_aib_txferclkoutn), .jtag_clkdr_in(clkdr_xr6r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp9),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_clkn), .oclkn(nc_oclkn_txferclkoutn),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top x446 ( .idata1_in1_jtag_out(idat1_poutp5),
     .async_dat_in1_jtag_out(nc_async_dat_poutp5),
     .idata0_in1_jtag_out(idat0_poutp5),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp5),
     .prev_io_shift_en(rshift_en_poutp[3]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_pout[5]), .oclk_out(nc_oclk[5]),
     .oclkb_out(nc_oclkb[5]), .odat0_out(nc_odat0[5]),
     .odat1_out(nc_odat1[5]), .odat_async_out(nc_odat_async[5]),
     .pd_data_out(nc_pd_data[5]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp5),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[5]),
     .idata0_in1(idat0_poutp3), .idata1_in0(idat1[5]),
     .idata1_in1(idat1_poutp3), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[0]), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk_r[2]),
     .ilaunch_clk_in1(tx_launch_clk_r[2]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp5), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[5]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[5]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_poutp5),
     .odat1_aib(nc_odat1_aib_pout[5]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp5),
     .odat0_aib(nc_odat0_aib_pout[5]), .oclk_aib(nc_oclk_aib_pout[5]),
     .last_bs_out(nc_last_bs_out_poutp5),
     .oclkb_aib(nc_oclkb_aib_pout[5]), .jtag_clkdr_in(clkdr_xr6r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp3),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[5]), .oclkn(nc_oclkn_pout[5]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top x438 ( .idata1_in1_jtag_out(idat1_poutp3),
     .async_dat_in1_jtag_out(nc_async_dat_poutp3),
     .idata0_in1_jtag_out(idat0_poutp3),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp3),
     .prev_io_shift_en(rshift_en_poutp[1]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_pout[3]), .oclk_out(nc_oclk[3]),
     .oclkb_out(nc_oclkb[3]), .odat0_out(nc_odat0[3]),
     .odat1_out(nc_odat1[3]), .odat_async_out(nc_odat_async[3]),
     .pd_data_out(nc_pd_data[3]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp3),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[3]),
     .idata0_in1(idat0_poutp1), .idata1_in0(idat1[3]),
     .idata1_in1(idat1_poutp1), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[0]), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk_r[6]),
     .ilaunch_clk_in1(tx_launch_clk_r[6]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp3), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[3]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[3]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_poutp3),
     .odat1_aib(nc_odat1_aib_pout[3]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp3),
     .odat0_aib(nc_odat0_aib_pout[3]), .oclk_aib(nc_oclk_aib_pout[3]),
     .last_bs_out(nc_last_bs_out_poutp3),
     .oclkb_aib(nc_oclkb_aib_pout[3]), .jtag_clkdr_in(clkdr_xr6r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp1),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[3]), .oclkn(nc_oclkn_pout[3]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top x430 ( .idata1_in1_jtag_out(idat1_poutp1),
     .async_dat_in1_jtag_out(nc_async_dat_poutp1),
     .idata0_in1_jtag_out(idat0_poutp1),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp1),
     .prev_io_shift_en(rshift_en_dtx[1]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(output_rstb), .pd_data_aib(nc_pd_data_aib_pout[1]),
     .oclk_out(nc_oclk[1]), .oclkb_out(nc_oclkb[1]),
     .odat0_out(nc_odat0[1]), .odat1_out(nc_odat1[1]),
     .odat_async_out(nc_odat_async[1]), .pd_data_out(nc_pd_data[1]),
     .async_dat_in0(vssl_aibnd), .async_dat_in1(async_dat_outpdir4_1),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp1),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[1]),
     .idata0_in1(vssl_aibnd), .idata1_in0(idat1[1]),
     .idata1_in1(vssl_aibnd), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[3]), .iddren_in0(iddren),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(tx_launch_clk_r[10]),
     .ilaunch_clk_in1(tx_launch_clk_r[10]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp1), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[3]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[1]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[1]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_poutp1),
     .odat1_aib(nc_odat1_aib_pout[1]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp1),
     .odat0_aib(nc_odat0_aib_pout[1]), .oclk_aib(nc_oclk_aib_pout[1]),
     .last_bs_out(nc_last_bs_out_poutp1),
     .oclkb_aib(nc_oclkb_aib_pout[1]), .jtag_clkdr_in(clkdr_xr6r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_outpdir4_1),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[1]), .oclkn(nc_oclkn_pout[1]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top x429 ( .idata1_in1_jtag_out(idat1_poutp7),
     .async_dat_in1_jtag_out(nc_async_dat_poutp7),
     .idata0_in1_jtag_out(idat0_poutp7),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp7),
     .prev_io_shift_en(rshift_en_poutp[5]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_pout[7]), .oclk_out(nc_oclk[7]),
     .oclkb_out(nc_oclkb[7]), .odat0_out(nc_odat0[7]),
     .odat1_out(nc_odat1[7]), .odat_async_out(nc_odat_async[7]),
     .pd_data_out(nc_pd_data[7]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp7),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[7]),
     .idata0_in1(idat0_poutp5), .idata1_in0(idat1[7]),
     .idata1_in1(idat1_poutp5), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[0]), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk_r[0]),
     .ilaunch_clk_in1(tx_launch_clk_r[0]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp7), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[7]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[7]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_poutp7),
     .odat1_aib(nc_odat1_aib_pout[7]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp7),
     .odat0_aib(nc_odat0_aib_pout[7]), .oclk_aib(nc_oclk_aib_pout[7]),
     .last_bs_out(nc_last_bs_out_poutp7),
     .oclkb_aib(nc_oclkb_aib_pout[7]), .jtag_clkdr_in(clkdr_xr6r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp5),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[7]), .oclkn(nc_oclkn_pout[7]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpoutp2 ( .idata1_in1_jtag_out(idat1_poutp2),
     .async_dat_in1_jtag_out(nc_async_dat_poutp2),
     .idata0_in1_jtag_out(idat0_poutp2),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp2),
     .prev_io_shift_en(rshift_en_poutp[0]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_pout[2]), .oclk_out(nc_oclk[2]),
     .oclkb_out(nc_oclkb[2]), .odat0_out(nc_odat0[2]),
     .odat1_out(nc_odat1[2]), .odat_async_out(nc_odat_async[2]),
     .pd_data_out(nc_pd_data[2]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp2),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[2]),
     .idata0_in1(idat0_poutp0), .idata1_in0(idat1[2]),
     .idata1_in1(idat1_poutp0), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[0]), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk_r[7]),
     .ilaunch_clk_in1(tx_launch_clk_r[7]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp2), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[2]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[2]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_poutp2),
     .odat1_aib(nc_odat1_aib_pout[2]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp2),
     .odat0_aib(nc_odat0_aib_pout[2]), .oclk_aib(nc_oclk_aib_pout[2]),
     .last_bs_out(nc_last_bs_out_poutp2),
     .oclkb_aib(nc_oclkb_aib_pout[2]), .jtag_clkdr_in(clkdr_xr5r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp0),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[2]), .oclkn(nc_oclkn_pout[2]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpoutp0 ( .idata1_in1_jtag_out(idat1_poutp0),
     .async_dat_in1_jtag_out(nc_async_dat_poutp0),
     .idata0_in1_jtag_out(idat0_poutp0),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp0),
     .prev_io_shift_en(shift_en_inpdir2), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(output_rstb), .pd_data_aib(nc_pd_data_aib_pout[0]),
     .oclk_out(nc_oclk[0]), .oclkb_out(nc_oclkb[0]),
     .odat0_out(nc_odat0[0]), .odat1_out(nc_odat1[0]),
     .odat_async_out(nc_odat_async[0]), .pd_data_out(nc_pd_data[0]),
     .async_dat_in0(vssl_aibnd), .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp0),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[0]),
     .idata0_in1(vssl_aibnd), .idata1_in0(idat1[0]),
     .idata1_in1(vssl_aibnd), .idataselb_in0(idataselb[0]),
     .idataselb_in1(vssl_aibnd), .iddren_in0(iddren),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(tx_launch_clk_r[11]),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1({vssl_aibnd, vssl_aibnd}), .irxen_in0({vssl_aibnd,
     vccl_aibnd, vssl_aibnd}), .irxen_in1(irxen_inpdir2[2:0]),
     .istrbclk_in0(jtag_clkdr_outn_poutp0), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(odat_async_pout0),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[0]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_poutp0),
     .odat1_aib(nc_odat1_aib_pout[0]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp0),
     .odat0_aib(nc_odat0_aib_pout[0]), .oclk_aib(nc_oclk_aib_pout[0]),
     .last_bs_out(nc_last_bs_out_poutp0),
     .oclkb_aib(nc_oclkb_aib_pout[0]), .jtag_clkdr_in(clkdr_xr5r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_directin2),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[0]), .oclkn(nc_oclkn_pout[0]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpoutp4 ( .idata1_in1_jtag_out(idat1_poutp4),
     .async_dat_in1_jtag_out(nc_async_dat_poutp4),
     .idata0_in1_jtag_out(idat0_poutp4),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp4),
     .prev_io_shift_en(rshift_en_poutp[2]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_pout[4]), .oclk_out(nc_oclk[4]),
     .oclkb_out(nc_oclkb[4]), .odat0_out(nc_odat0[4]),
     .odat1_out(nc_odat1[4]), .odat_async_out(nc_odat_async[4]),
     .pd_data_out(nc_pd_data[4]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp4),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[4]),
     .idata0_in1(idat0_poutp2), .idata1_in0(idat1[4]),
     .idata1_in1(idat1_poutp2), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[0]), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk_r[3]),
     .ilaunch_clk_in1(tx_launch_clk_r[3]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp4), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[4]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[4]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_poutp4),
     .odat1_aib(nc_odat1_aib_pout[4]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp4),
     .odat0_aib(nc_odat0_aib_pout[4]), .oclk_aib(nc_oclk_aib_pout[4]),
     .last_bs_out(nc_last_bs_out_poutp4),
     .oclkb_aib(nc_oclkb_aib_pout[4]), .jtag_clkdr_in(clkdr_xr5r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp2),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[4]), .oclkn(nc_oclkn_pout[4]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpoutp11 ( .idata1_in1_jtag_out(idat1_poutp11),
     .async_dat_in1_jtag_out(nc_async_dat_poutp11),
     .idata0_in1_jtag_out(idat0_poutp11),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp11),
     .prev_io_shift_en(rshift_en_txferclkoutn),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_pout[11]), .oclk_out(nc_oclk[11]),
     .oclkb_out(nc_oclkb[11]), .odat0_out(nc_odat0[11]),
     .odat1_out(nc_odat1[11]), .odat_async_out(nc_odat_async[11]),
     .pd_data_out(nc_pd_data[11]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp11),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[11]),
     .idata0_in1(idata0_in1_clkn), .idata1_in0(idat1[11]),
     .idata1_in1(idata1_in1_clkn), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[1]), .iddren_in0(iddren),
     .iddren_in1(vccl_aibnd), .ilaunch_clk_in0(tx_launch_clk_l[10]),
     .ilaunch_clk_in1(tx_launch_clk_l[10]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp11), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[1]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[11]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[11]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_poutp11),
     .odat1_aib(nc_odat1_aib_pout[11]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp11),
     .odat0_aib(nc_odat0_aib_pout[11]),
     .oclk_aib(nc_oclk_aib_pout[11]),
     .last_bs_out(nc_last_bs_out_poutp11),
     .oclkb_aib(nc_oclkb_aib_pout[11]), .jtag_clkdr_in(clkdr_xr6l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_clkn),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[11]), .oclkn(nc_oclkn_pout[11]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xasyncrx0 ( .idata1_in1_jtag_out(nc_idat1_inpshared0),
     .async_dat_in1_jtag_out(nc_async_dat_inpshared0),
     .idata0_in1_jtag_out(nc_idat0_inpshared0),
     .jtag_clkdr_outn(jtag_clkdr_outn_inpshared0),
     .prev_io_shift_en(rshift_en_tx[2]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(output_rstb), .pd_data_aib(ncrx_pd_data_aib[0]),
     .oclk_out(odat_async[0]), .oclkb_out(ncrx_oclkb[0]),
     .odat0_out(ncrx_odat0[0]), .odat1_out(ncrx_odat1[0]),
     .odat_async_out(ncrx_async_data_out0),
     .pd_data_out(ncrx_pd_data[0]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(vssl_aibnd),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vssl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(oclk_inpdir2), .odat_async_aib(ncrx_odat_async_aib[0]),
     .oclkb_in1(oclkb_inpdir2), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_tx[0]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(output_rstb), .jtag_clkdr_out(jtag_clkdr_inpshared0),
     .odat1_aib(ncrx_odat1_aib[0]),
     .jtag_rx_scan_out(jtag_rx_scan_inpshared0),
     .odat0_aib(ncrx_odat0_aib[0]), .oclk_aib(oclk_inpshared0),
     .last_bs_out(nc_last_bs_out_diro0), .oclkb_aib(oclkb_inpshared0),
     .jtag_clkdr_in(clkdr_xr3r), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_async_in2),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_async_in[0]), .oclkn(ncrx_oclkn0),
     .iclkn(oclkn_inpshared1), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdirect_in2 ( .idata1_in1_jtag_out(nc_idat1_inpclk3),
     .async_dat_in1_jtag_out(nc_async_dat_inpclk3),
     .idata0_in1_jtag_out(nc_idat0_inpclk3),
     .jtag_clkdr_outn(jtag_clkdr_outn_inpclk3),
     .prev_io_shift_en(shift_en_inpclk1n), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(output_rstb), .pd_data_aib(ncdrx_pd_data_aib[2]),
     .oclk_out(ncdrx_oclk[2]), .oclkb_out(ncdrx_oclkb[2]),
     .odat0_out(ncdrx_odat0[2]), .odat1_out(ncdrx_odat1[2]),
     .odat_async_out(odirectin_data[2]),
     .pd_data_out(ncdrx_pd_data[2]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(vssl_aibnd),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vssl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r1[2:0]), .irxen_in1({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .istrbclk_in0(vssl_aibnd),
     .istrbclk_in1(vssl_aibnd), .itxen_in0(vssl_aibnd),
     .itxen_in1(vssl_aibnd), .oclk_in1(vssl_aibnd),
     .odat_async_aib(ncdrx_odat_async_aib[2]), .oclkb_in1(vssl_aibnd),
     .odat0_in1(vssl_aibnd), .odat1_in1(vssl_aibnd),
     .odat_async_in1(odat_async_inpclk4), .shift_en(rshift_en_drx[2]),
     .pd_data_in1(vssl_aibnd), .dig_rstb(output_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_inpclk3),
     .odat1_aib(ncdrx_odat1_aib[2]),
     .jtag_rx_scan_out(jtag_rx_scan_out_inpclk3),
     .odat0_aib(ncdrx_odat0_aib2), .oclk_aib(oclk_inpclk3),
     .last_bs_out(nc_last_bs_out_inpclk3), .oclkb_aib(oclkb_inpclk3),
     .jtag_clkdr_in(clkdr_xr2l), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_inpclk1n),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_direct_input[2]), .oclkn(oclkn_inpclk3),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdirect_out3 (
     .idata1_in1_jtag_out(nc_idat1_outpdir1_1),
     .async_dat_in1_jtag_out(async_dat_outpdir1_1),
     .idata0_in1_jtag_out(nc_idat0_outpdir1_1),
     .jtag_clkdr_outn(jtag_clkdr_outn_outpdir1_1),
     .prev_io_shift_en(shift_en_outpclk0), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(output_rstb), .pd_data_aib(ncdtx_pd_data_aib[3]),
     .oclk_out(ncdtx_oclk[3]), .oclkb_out(ncdtx_oclkb[3]),
     .odat0_out(ncdtx_odat0[3]), .odat1_out(ncdtx_odat1[3]),
     .odat_async_out(ncdtx_odat_async[3]),
     .pd_data_out(ncdtx_pd_data[3]),
     .async_dat_in0(idirectout_data[3]), .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(vssl_aibnd), .iclkin_dist_in1(vssl_aibnd),
     .idata0_in0(vssl_aibnd), .idata0_in1(idat0_in0_dout_clkp),
     .idata1_in0(vssl_aibnd), .idata1_in1(idat1_in0_dout_clkp),
     .idataselb_in0(idataselb[3]),
     .idataselb_in1(idataselb_in0_dout_clkp), .iddren_in0(vssl_aibnd),
     .iddren_in1(vccl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(ilaunch_clk_in0_dout_clkp),
     .ilpbk_dat_in0(vssl_aibnd), .ilpbk_dat_in1(vssl_aibnd),
     .ilpbk_en_in0(vssl_aibnd), .ilpbk_en_in1(vssl_aibnd),
     .indrv_in0(indrv_r34[1:0]), .indrv_in1(indrv_r34[1:0]),
     .ipdrv_in0(ipdrv_r34[1:0]), .ipdrv_in1(ipdrv_r34[1:0]),
     .irxen_in0({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[3]), .itxen_in1(itxen_in0_dout_clkp),
     .oclk_in1(vssl_aibnd), .odat_async_aib(ncdtx_odat_async_aib3),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_dtx[3]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(output_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_outpdir1_1),
     .odat1_aib(ncdtx_odat1_aib[3]),
     .jtag_rx_scan_out(jtag_rx_scan_out_outpdir1_1),
     .odat0_aib(ncdtx_odat0_aib[3]), .oclk_aib(ncdtx_oclk_aib[3]),
     .last_bs_out(nc_last_bs_out_outpdir1_1),
     .oclkb_aib(ncdtx_oclkb_aib3), .jtag_clkdr_in(clkdr_xr3l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_diin_clkp),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_directout[3]), .oclkn(ncdtx_oclkn[3]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpoutp6 ( .idata1_in1_jtag_out(idat1_poutp6),
     .async_dat_in1_jtag_out(nc_async_dat_poutp6),
     .idata0_in1_jtag_out(idat0_poutp6),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp6),
     .prev_io_shift_en(rshift_en_poutp[4]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_pout[6]), .oclk_out(nc_oclk[6]),
     .oclkb_out(nc_oclkb[6]), .odat0_out(nc_odat0[6]),
     .odat1_out(nc_odat1[6]), .odat_async_out(nc_odat_async[6]),
     .pd_data_out(nc_pd_data[6]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp6),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[6]),
     .idata0_in1(idat0_poutp4), .idata1_in0(idat1[6]),
     .idata1_in1(idat1_poutp4), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[0]), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk_r[1]),
     .ilaunch_clk_in1(tx_launch_clk_r[1]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp6), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[6]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[6]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_poutp6),
     .odat1_aib(nc_odat1_aib_pout[6]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp6),
     .odat0_aib(nc_odat0_aib_pout[6]), .oclk_aib(nc_oclk_aib_pout[6]),
     .last_bs_out(nc_last_bs_out_poutp6),
     .oclkb_aib(nc_oclkb_aib_pout[6]), .jtag_clkdr_in(clkdr_xr5r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp4),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[6]), .oclkn(nc_oclkn_pout[6]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpoutp8 ( .idata1_in1_jtag_out(idat1_poutp8),
     .async_dat_in1_jtag_out(nc_async_dat_poutp8),
     .idata0_in1_jtag_out(idat0_poutp8),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp8),
     .prev_io_shift_en(rshift_en_poutp[6]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_pout[8]), .oclk_out(nc_oclk[8]),
     .oclkb_out(nc_oclkb[8]), .odat0_out(nc_odat0[8]),
     .odat1_out(nc_odat1[8]), .odat_async_out(nc_odat_async[8]),
     .pd_data_out(nc_pd_data[8]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp8),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[8]),
     .idata0_in1(idat0_poutp6), .idata1_in0(idat1[8]),
     .idata1_in1(idat1_poutp6), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[0]), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk_r[5]),
     .ilaunch_clk_in1(tx_launch_clk_r[5]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp8), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[8]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[8]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_poutp8),
     .odat1_aib(nc_odat1_aib_pout[8]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp8),
     .odat0_aib(nc_odat0_aib_pout[8]), .oclk_aib(nc_oclk_aib_pout[8]),
     .last_bs_out(nc_last_bs_out_poutp8),
     .oclkb_aib(nc_oclkb_aib_pout[8]), .jtag_clkdr_in(clkdr_xr5r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp6),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[8]), .oclkn(nc_oclkn_pout[8]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top x187 ( .idata1_in1_jtag_out(idata1_in1_clkp),
     .async_dat_in1_jtag_out(nc_async_dat_clkp),
     .idata0_in1_jtag_out(idata0_in1_clkp),
     .jtag_clkdr_outn(jtag_clkdr_outn_clkp),
     .prev_io_shift_en(rshift_en_poutp[8]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_txferclkout), .oclk_out(nc_oclk_clkp),
     .oclkb_out(nc_oclkb_clkp), .odat0_out(nc_odat0_clkp),
     .odat1_out(nc_odat1_clkp), .odat_async_out(nc_odat_async_clkp),
     .pd_data_out(nc_pd_data_clkp), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_clkp),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0_clkp),
     .idata0_in1(idat0_poutp8), .idata1_in0(idat1_clkp),
     .idata1_in1(idat1_poutp8), .idataselb_in0(idataselb[1]),
     .idataselb_in1(idataselb[0]), .iddren_in0(vccl_aibnd),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk_r[9]),
     .ilaunch_clk_in1(tx_launch_clk_r[9]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_clkp), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[1]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_txferclkout),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_txferclkout), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_clkp),
     .odat1_aib(nc_odat1_aib_txferclkout),
     .jtag_rx_scan_out(jtag_rx_scan_out_clkp),
     .odat0_aib(nc_odat0_aib_txferclkout),
     .oclk_aib(nc_oclk_aib_txferclkout),
     .last_bs_out(nc_last_bs_out_txferclkout),
     .oclkb_aib(nc_oclkb_aib_txferclkout), .jtag_clkdr_in(clkdr_xr5r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp8),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_clkp), .oclkn(nc_oclkn_txferclkout),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpoutp10 ( .idata1_in1_jtag_out(idat1_poutp10),
     .async_dat_in1_jtag_out(nc_async_dat_poutp10),
     .idata0_in1_jtag_out(idat0_poutp10),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp10),
     .prev_io_shift_en(rshift_en_txferclkout),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_pout[10]), .oclk_out(nc_oclk[10]),
     .oclkb_out(nc_oclkb[10]), .odat0_out(nc_odat0[10]),
     .odat1_out(nc_odat1[10]), .odat_async_out(nc_odat_async[10]),
     .pd_data_out(nc_pd_data[10]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp10),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[10]),
     .idata0_in1(idata0_in1_clkp), .idata1_in0(idat1[10]),
     .idata1_in1(idata1_in1_clkp), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[1]), .iddren_in0(iddren),
     .iddren_in1(vccl_aibnd), .ilaunch_clk_in0(tx_launch_clk_l[11]),
     .ilaunch_clk_in1(tx_launch_clk_l[11]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp10), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[1]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[10]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[10]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_poutp10),
     .odat1_aib(nc_odat1_aib_pout[10]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp10),
     .odat0_aib(nc_odat0_aib_pout[10]),
     .oclk_aib(nc_oclk_aib_pout[10]),
     .last_bs_out(nc_last_bs_out_poutp10),
     .oclkb_aib(nc_oclkb_aib_pout[10]), .jtag_clkdr_in(clkdr_xr5l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_clkp),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[10]), .oclkn(nc_oclkn_pout[10]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpoutp12 ( .idata1_in1_jtag_out(idat1_poutp12),
     .async_dat_in1_jtag_out(nc_async_dat_poutp12),
     .idata0_in1_jtag_out(idat0_poutp12),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp12),
     .prev_io_shift_en(rshift_en_poutp[10]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_pout[12]), .oclk_out(nc_oclk[12]),
     .oclkb_out(nc_oclkb[12]), .odat0_out(nc_odat0[12]),
     .odat1_out(nc_odat1[12]), .odat_async_out(nc_odat_async[12]),
     .pd_data_out(nc_pd_data[12]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp12),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[12]),
     .idata0_in1(idat0_poutp10), .idata1_in0(idat1[12]),
     .idata1_in1(idat1_poutp10), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[0]), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk_l[7]),
     .ilaunch_clk_in1(tx_launch_clk_l[7]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp12), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[12]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[12]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_poutp12),
     .odat1_aib(nc_odat1_aib_pout[12]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp12),
     .odat0_aib(nc_odat0_aib_pout[12]),
     .oclk_aib(nc_oclk_aib_pout[12]),
     .last_bs_out(nc_last_bs_out_poutp12),
     .oclkb_aib(nc_oclkb_aib_pout[12]), .jtag_clkdr_in(clkdr_xr5l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp10),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[12]), .oclkn(nc_oclkn_pout[12]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpoutp13 ( .idata1_in1_jtag_out(idat1_poutp13),
     .async_dat_in1_jtag_out(nc_async_dat_poutp13),
     .idata0_in1_jtag_out(idat0_poutp13),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp13),
     .prev_io_shift_en(rshift_en_poutp[11]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_pout[13]), .oclk_out(nc_oclk[13]),
     .oclkb_out(nc_oclkb[13]), .odat0_out(nc_odat0[13]),
     .odat1_out(nc_odat1[13]), .odat_async_out(nc_odat_async[13]),
     .pd_data_out(nc_pd_data[13]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp13),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[13]),
     .idata0_in1(idat0_poutp11), .idata1_in0(idat1[13]),
     .idata1_in1(idat1_poutp11), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[0]), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk_l[6]),
     .ilaunch_clk_in1(tx_launch_clk_l[6]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp13), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[13]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[13]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_poutp13),
     .odat1_aib(nc_odat1_aib_pout[13]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp13),
     .odat0_aib(nc_odat0_aib_pout[13]),
     .oclk_aib(nc_oclk_aib_pout[13]),
     .last_bs_out(nc_last_bs_out_poutp13),
     .oclkb_aib(nc_oclkb_aib_pout[13]), .jtag_clkdr_in(clkdr_xr6l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp11),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[13]), .oclkn(nc_oclkn_pout[13]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpoutp14 ( .idata1_in1_jtag_out(idat1_poutp14),
     .async_dat_in1_jtag_out(nc_async_dat_poutp14),
     .idata0_in1_jtag_out(idat0_poutp14),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp14),
     .prev_io_shift_en(rshift_en_poutp[12]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_pout[14]), .oclk_out(nc_oclk[14]),
     .oclkb_out(nc_oclkb[14]), .odat0_out(nc_odat0[14]),
     .odat1_out(nc_odat1[14]), .odat_async_out(nc_odat_async[14]),
     .pd_data_out(nc_pd_data[14]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp14),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[14]),
     .idata0_in1(idat0_poutp12), .idata1_in0(idat1[14]),
     .idata1_in1(idat1_poutp12), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[0]), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk_l[3]),
     .ilaunch_clk_in1(tx_launch_clk_l[3]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp14), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[14]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[14]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_poutp14),
     .odat1_aib(nc_odat1_aib_pout[14]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp14),
     .odat0_aib(nc_odat0_aib_pout[14]),
     .oclk_aib(nc_oclk_aib_pout[14]),
     .last_bs_out(nc_last_bs_out_poutp14),
     .oclkb_aib(nc_oclkb_aib_pout[14]), .jtag_clkdr_in(clkdr_xr5l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp12),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[14]), .oclkn(nc_oclkn_pout[14]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpoutp15 ( .idata1_in1_jtag_out(idat1_poutp15),
     .async_dat_in1_jtag_out(nc_async_dat_poutp15),
     .idata0_in1_jtag_out(idat0_poutp15),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp15),
     .prev_io_shift_en(rshift_en_poutp[13]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_pout[15]), .oclk_out(nc_oclk[15]),
     .oclkb_out(nc_oclkb[15]), .odat0_out(nc_odat0[15]),
     .odat1_out(nc_odat1[15]), .odat_async_out(nc_odat_async[15]),
     .pd_data_out(nc_pd_data[15]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp15),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[15]),
     .idata0_in1(idat0_poutp13), .idata1_in0(idat1[15]),
     .idata1_in1(idat1_poutp13), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[0]), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk_l[2]),
     .ilaunch_clk_in1(tx_launch_clk_l[2]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp15), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[15]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[15]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_poutp15),
     .odat1_aib(nc_odat1_aib_pout[15]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp15),
     .odat0_aib(nc_odat0_aib_pout[15]),
     .oclk_aib(nc_oclk_aib_pout[15]),
     .last_bs_out(nc_last_bs_out_poutp15),
     .oclkb_aib(nc_oclkb_aib_pout[15]), .jtag_clkdr_in(clkdr_xr6l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp13),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[15]), .oclkn(nc_oclkn_pout[15]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdirect_in0 ( .idata1_in1_jtag_out(nc_idat1_inpdir3),
     .async_dat_in1_jtag_out(nc_async_dat_inpdir3),
     .idata0_in1_jtag_out(nc_idat0_inpdir3),
     .jtag_clkdr_outn(jtag_clkdr_outn_inpdir3),
     .prev_io_shift_en(rshift_en_dirclkp[1]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(ncdrx_pd_data_aib[0]), .oclk_out(ncdrx_oclk[0]),
     .oclkb_out(ncdrx_oclkb[0]), .odat0_out(ncdrx_odat0[0]),
     .odat1_out(ncdrx_odat1[0]), .odat_async_out(odirectin_data[0]),
     .pd_data_out(ncdrx_pd_data[0]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(vssl_aibnd),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vssl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r1[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(ncdrx_odat_async_aib[0]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(odat_async_inpclk1),
     .shift_en(rshift_en_drx[0]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(output_rstb), .jtag_clkdr_out(jtag_clkdr_out_inpdir3),
     .odat1_aib(ncdrx_odat1_aib0),
     .jtag_rx_scan_out(jtag_rx_scan_out_inpdir3),
     .odat0_aib(ncdrx_odat0_aib[0]), .oclk_aib(drx_oclk_aib[0]),
     .last_bs_out(nc_last_bs_out_inpdir3),
     .oclkb_aib(drx_oclkb_aib[0]), .jtag_clkdr_in(clkdr_xr1l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_dirclkp1),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_direct_input[0]), .oclkn(ncdrx_oclkn0),
     .iclkn(oclkn_inpdir4), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xasynctx1 ( .idata1_in1_jtag_out(nc_idat1_async_out1),
     .async_dat_in1_jtag_out(async_dat_async_out1),
     .idata0_in1_jtag_out(nc_idat0_async_out1),
     .jtag_clkdr_outn(jtag_clkdr_outn_async_out1),
     .prev_io_shift_en(shift_en_inpclk6), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(output_rstb), .pd_data_aib(nctx_pd_data_aib[1]),
     .oclk_out(nctx_oclk[1]), .oclkb_out(nctx_oclkb[1]),
     .odat0_out(nctx_odat0[1]), .odat1_out(nctx_odat1[1]),
     .odat_async_out(nctx_odat_async[1]),
     .pd_data_out(nctx_pd_data[1]), .async_dat_in0(iasyncdata[1]),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(vssl_aibnd),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(idataselb[2]),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r12[1:0]),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0(ipdrv_r12[1:0]),
     .ipdrv_in1({vssl_aibnd, vssl_aibnd}), .irxen_in0({vssl_aibnd,
     vccl_aibnd, vssl_aibnd}), .irxen_in1(irxen_inpclk6[2:0]),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[2]), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(odat_async_oshared1),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(odat_async_aib2),
     .shift_en(rshift_en_rx[1]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(output_rstb), .jtag_clkdr_out(jtag_clkdr_async_out1),
     .odat1_aib(nctx_odat1_aib[1]),
     .jtag_rx_scan_out(jtag_rx_scan_async_out1),
     .odat0_aib(nctx_odat0_aib[1]), .oclk_aib(nctx_oclk_aib[1]),
     .last_bs_out(nc_last_bs_out_oshared1),
     .oclkb_aib(nctx_oclkb_aib[1]), .jtag_clkdr_in(clkdr_xr2r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_inpclk6),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_async_out[1]), .oclkn(nctx_oclkn[1]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xasynctx2 ( .idata1_in1_jtag_out(nc_idat1_async_out2),
     .async_dat_in1_jtag_out(iasyncdata_oshared2),
     .idata0_in1_jtag_out(nc_idat0_async_out2),
     .jtag_clkdr_outn(jtag_clkdr_outn_async_out2),
     .prev_io_shift_en(rshift_en_rx[1]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(output_rstb), .pd_data_aib(nctx_pd_data_aib[2]),
     .oclk_out(nctx_oclk[2]), .oclkb_out(nctx_oclkb[2]),
     .odat0_out(nctx_odat0[2]), .odat1_out(nctx_odat1[2]),
     .odat_async_out(nctx_odat_async[2]),
     .pd_data_out(nctx_pd_data[2]), .async_dat_in0(iasyncdata[2]),
     .async_dat_in1(async_dat_async_out1),
     .iclkin_dist_in0(vssl_aibnd), .iclkin_dist_in1(vssl_aibnd),
     .idata0_in0(vssl_aibnd), .idata0_in1(vssl_aibnd),
     .idata1_in0(vssl_aibnd), .idata1_in1(vssl_aibnd),
     .idataselb_in0(idataselb[2]), .idataselb_in1(idataselb[2]),
     .iddren_in0(vssl_aibnd), .iddren_in1(vssl_aibnd),
     .ilaunch_clk_in0(vssl_aibnd), .ilaunch_clk_in1(vssl_aibnd),
     .ilpbk_dat_in0(vssl_aibnd), .ilpbk_dat_in1(vssl_aibnd),
     .ilpbk_en_in0(vssl_aibnd), .ilpbk_en_in1(vssl_aibnd),
     .indrv_in0(indrv_r12[1:0]), .indrv_in1(indrv_r12[1:0]),
     .ipdrv_in0(ipdrv_r12[1:0]), .ipdrv_in1(ipdrv_r12[1:0]),
     .irxen_in0({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[2]), .itxen_in1(itxen[2]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(odat_async_aib2), .oclkb_in1(vssl_aibnd),
     .odat0_in1(vssl_aibnd), .odat1_in1(vssl_aibnd),
     .odat_async_in1(vssl_aibnd), .shift_en(rshift_en_rx[3]),
     .pd_data_in1(vssl_aibnd), .dig_rstb(output_rstb),
     .jtag_clkdr_out(jtag_clkdr_oshared2),
     .odat1_aib(nctx_odat1_aib[2]),
     .jtag_rx_scan_out(jtag_rx_scan_oshared2),
     .odat0_aib(nctx_odat0_aib[2]), .oclk_aib(nctx_oclk_aib[2]),
     .last_bs_out(nc_last_bs_out_oshared2),
     .oclkb_aib(nctx_oclkb_aib[2]), .jtag_clkdr_in(clkdr_xr2r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_async_out1),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_async_out[2]), .oclkn(nctx_oclkn[2]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xasyncrx4 ( .idata1_in1_jtag_out(nc_idat1_inpshared4),
     .async_dat_in1_jtag_out(nc_async_dat_inpshared4),
     .idata0_in1_jtag_out(nc_idat0_inpshared4),
     .jtag_clkdr_outn(jtag_clkdr_outn_inpshared4),
     .prev_io_shift_en(rshift_en_rx[0]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(output_rstb), .pd_data_aib(ncrx_pd_data_aib[4]),
     .oclk_out(ncrx_oclk[4]), .oclkb_out(ncrx_oclkb[4]),
     .odat0_out(ncrx_odat0[4]), .odat1_out(ncrx_odat1[4]),
     .odat_async_out(odat_async[4]), .pd_data_out(ncrx_pd_data[4]),
     .async_dat_in0(vssl_aibnd), .async_dat_in1(async_dat_async_out0),
     .iclkin_dist_in0(vssl_aibnd), .iclkin_dist_in1(vssl_aibnd),
     .idata0_in0(vssl_aibnd), .idata0_in1(vssl_aibnd),
     .idata1_in0(vssl_aibnd), .idata1_in1(vssl_aibnd),
     .idataselb_in0(vssl_aibnd), .idataselb_in1(idataselb[2]),
     .iddren_in0(vssl_aibnd), .iddren_in1(vssl_aibnd),
     .ilaunch_clk_in0(vssl_aibnd), .ilaunch_clk_in1(vssl_aibnd),
     .ilpbk_dat_in0(vssl_aibnd), .ilpbk_dat_in1(vssl_aibnd),
     .ilpbk_en_in0(vssl_aibnd), .ilpbk_en_in1(vssl_aibnd),
     .indrv_in0({vssl_aibnd, vssl_aibnd}), .indrv_in1(indrv_r12[1:0]),
     .ipdrv_in0({vssl_aibnd, vssl_aibnd}), .ipdrv_in1(ipdrv_r12[1:0]),
     .irxen_in0(irxen_r2[2:0]), .irxen_in1({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .istrbclk_in0(vssl_aibnd),
     .istrbclk_in1(vssl_aibnd), .itxen_in0(vssl_aibnd),
     .itxen_in1(itxen[2]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(odat_async_aib4), .oclkb_in1(vssl_aibnd),
     .odat0_in1(vssl_aibnd), .odat1_in1(vssl_aibnd),
     .odat_async_in1(odat_async_fsrdin), .shift_en(rshift_en_rx[2]),
     .pd_data_in1(vssl_aibnd), .dig_rstb(output_rstb),
     .jtag_clkdr_out(jtag_clkdr_inpshared4),
     .odat1_aib(ncrx_odat1_aib[4]),
     .jtag_rx_scan_out(jtag_rx_scan_inpshared4),
     .odat0_aib(ncrx_odat0_aib[4]), .oclk_aib(ncrx_oclk_aib[4]),
     .last_bs_out(nc_last_bs_out_inpshared4),
     .oclkb_aib(ncrx_oclkb_aib[4]), .jtag_clkdr_in(clkdr_xr1r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_async_out0),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_async_in[4]), .oclkn(ncrx_oclkn4),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top x740 ( .idata1_in1_jtag_out(nc_idat1_ptxclkinn),
     .async_dat_in1_jtag_out(nc_async_dat_ptxclkinn),
     .idata0_in1_jtag_out(nc_idat0_ptxclkinn),
     .jtag_clkdr_outn(jtag_clkdr_outn_ptxclkinn),
     .prev_io_shift_en(shift_en_voutp01), .anlg_rstb(output_rstb),
     .pd_data_aib(ncrx_pd_data_aib_clkn0),
     .oclk_out(ncout_rx_fast_clkn[0]),
     .oclkb_out(ncout_rx_fast_clknb[0]),
     .odat0_out(nc_rxodat0_clkn[0]), .odat1_out(nc_rxodat1_clkn[0]),
     .odat_async_out(nc_rxodat_async_clkn[0]),
     .pd_data_out(nc_rxpd_data_clkn[0]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(vssl_aibnd),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(idat0_voutp01), .idata1_in0(vssl_aibnd),
     .idata1_in1(idat1_voutp01), .idataselb_in0(vssl_aibnd),
     .idataselb_in1(idataselb_voutp01), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(ilaunch_clk_voutp01), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1(indrv_r34[1:0]), .ipdrv_in0({vssl_aibnd, vssl_aibnd}),
     .ipdrv_in1(ipdrv_r34[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(vssl_aibnd), .itxen_in1(itxen_voutp01),
     .oclk_in1(vssl_aibnd), .odat_async_aib(ncrx_odat_async_aib_clkn0),
     .oclkb_in1(vssl_aibnd), .jtag_clksel(jtag_clksel),
     .odat0_in1(vssl_aibnd), .vssl_aibnd(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_dirclkn[0]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(avmm_sync_rstb), .jtag_clkdr_out(jtag_clkdr_ptxclkinn),
     .jtag_intest(jtag_intest), .odat1_aib(ncrx_odat1_aib_clkn0),
     .jtag_rx_scan_out(jtag_rx_scan_ptxclkinn),
     .odat0_aib(ncrx_odat0_aib_clkn0),
     .oclk_aib(nc_out_rx_fast_clkn_aib0),
     .last_bs_out(nc_last_bs_out_ptxclkinn), .vccl_aibnd(vccl_aibnd),
     .oclkb_aib(nc_out_rx_fast_clknb_aib0), .jtag_clkdr_in(clkdr_xr4l),
     .jtag_rstb_en(jtag_rstb_en), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_voutp01),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_directinclkn[0]), .oclkn(oclkn_clkn0),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdirect_out1 (
     .idata1_in1_jtag_out(nc_idat1_outpdir4_1),
     .async_dat_in1_jtag_out(async_dat_outpdir4_1),
     .idata0_in1_jtag_out(nc_idat0_outpdir4_1),
     .jtag_clkdr_outn(jtag_clkdr_outn_outpdir4_1),
     .prev_io_shift_en(rshift_en_tx[1]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(output_rstb), .pd_data_aib(ncdtx_pd_data_aib[1]),
     .oclk_out(ncdtx_oclk[1]), .oclkb_out(ncdtx_oclkb[1]),
     .odat0_out(ncdtx_odat0[1]), .odat1_out(ncdtx_odat1[1]),
     .odat_async_out(ncdtx_odat_async[1]),
     .pd_data_out(ncdtx_pd_data[1]),
     .async_dat_in0(idirectout_data[1]), .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(vssl_aibnd), .iclkin_dist_in1(vssl_aibnd),
     .idata0_in0(vssl_aibnd), .idata0_in1(vssl_aibnd),
     .idata1_in0(vssl_aibnd), .idata1_in1(vssl_aibnd),
     .idataselb_in0(idataselb[3]), .idataselb_in1(vssl_aibnd),
     .iddren_in0(vssl_aibnd), .iddren_in1(vssl_aibnd),
     .ilaunch_clk_in0(vssl_aibnd), .ilaunch_clk_in1(vssl_aibnd),
     .ilpbk_dat_in0(vssl_aibnd), .ilpbk_dat_in1(vssl_aibnd),
     .ilpbk_en_in0(vssl_aibnd), .ilpbk_en_in1(vssl_aibnd),
     .indrv_in0(indrv_r34[1:0]), .indrv_in1({vssl_aibnd, vssl_aibnd}),
     .ipdrv_in0(ipdrv_r34[1:0]), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[3]), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(ncdtx_odat_async_aib[1]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_dtx[1]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(output_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_outpdir4_1),
     .odat1_aib(ncdtx_odat1_aib[1]),
     .jtag_rx_scan_out(jtag_rx_scan_out_outpdir4_1),
     .odat0_aib(ncdtx_odat0_aib[1]), .oclk_aib(ncdtx_oclk_aib1),
     .last_bs_out(nc_last_bs_out_outpdir4_1),
     .oclkb_aib(ncdtx_oclkb_aib[1]), .jtag_clkdr_in(clkdr_xr4r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_async_in1),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_directout[1]), .oclkn(dtx_oclkn1),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpoutp18 ( .idata1_in1_jtag_out(idat1_poutp18),
     .async_dat_in1_jtag_out(nc_async_dat_poutp18),
     .idata0_in1_jtag_out(idat0_poutp18),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp18),
     .prev_io_shift_en(rshift_en_poutp[16]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_pout[18]), .oclk_out(nc_oclk[18]),
     .oclkb_out(nc_oclkb[18]), .odat0_out(nc_odat0[18]),
     .odat1_out(nc_odat1[18]), .odat_async_out(nc_odat_async[18]),
     .pd_data_out(nc_pd_data[18]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp18),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[18]),
     .idata0_in1(idat0_poutp16), .idata1_in0(idat1[18]),
     .idata1_in1(idat1_poutp16), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[0]), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk_l[5]),
     .ilaunch_clk_in1(tx_launch_clk_l[5]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp18), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[18]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[18]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_poutp18),
     .odat1_aib(nc_odat1_aib_pout[18]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp18),
     .odat0_aib(nc_odat0_aib_pout[18]),
     .oclk_aib(nc_oclk_aib_pout[18]),
     .last_bs_out(nc_last_bs_out_poutp18),
     .oclkb_aib(nc_oclkb_aib_pout[18]), .jtag_clkdr_in(clkdr_xr5l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp16),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[18]), .oclkn(nc_oclkn_pout[18]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdiin_clkn ( .idata1_in1_jtag_out(nc_idat1_inpclk0n),
     .async_dat_in1_jtag_out(nc_async_dat_inpclk0n),
     .idata0_in1_jtag_out(nc_idat0_inpclk0n),
     .jtag_clkdr_outn(jtag_clkdr_outn_inpclk0n),
     .prev_io_shift_en(shift_en_outpdir0_1),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(ncrx_pd_data_aib_clkn1),
     .oclk_out(ncout_rx_fast_clkn[1]),
     .oclkb_out(ncout_rx_fast_clknb[1]),
     .odat0_out(nc_rxodat0_clkn[1]), .odat1_out(nc_rxodat1_clkn[1]),
     .odat_async_out(nc_rxodat_async_clkn[1]),
     .pd_data_out(nc_rxpd_data_clkn[1]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(async_dat_outpdir0_1),
     .iclkin_dist_in0(vssl_aibnd), .iclkin_dist_in1(vssl_aibnd),
     .idata0_in0(vssl_aibnd), .idata0_in1(vssl_aibnd),
     .idata1_in0(vssl_aibnd), .idata1_in1(vssl_aibnd),
     .idataselb_in0(vssl_aibnd), .idataselb_in1(idataselb_outpdir0_1),
     .iddren_in0(vssl_aibnd), .iddren_in1(vssl_aibnd),
     .ilaunch_clk_in0(vssl_aibnd), .ilaunch_clk_in1(vssl_aibnd),
     .ilpbk_dat_in0(vssl_aibnd), .ilpbk_dat_in1(vssl_aibnd),
     .ilpbk_en_in0(vssl_aibnd), .ilpbk_en_in1(vssl_aibnd),
     .indrv_in0({vssl_aibnd, vssl_aibnd}), .indrv_in1(indrv_r12[1:0]),
     .ipdrv_in0({vssl_aibnd, vssl_aibnd}), .ipdrv_in1(ipdrv_r12[1:0]),
     .irxen_in0({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(vssl_aibnd), .itxen_in1(itxen_outpdir0_1),
     .oclk_in1(vssl_aibnd), .odat_async_aib(ncrx_odat_async_aib_clkn1),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_dirclkn[1]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(output_rstb), .jtag_clkdr_out(jtag_clkdr_inpclk0n),
     .odat1_aib(ncrx_odat1_aib_clkn1),
     .jtag_rx_scan_out(jtag_rx_scan_inpclk0n),
     .odat0_aib(ncrx_odat0_aib_clkn1),
     .oclk_aib(nc_out_rx_fast_clkn_aib1),
     .last_bs_out(nc_last_bs_out_inpclk0n),
     .oclkb_aib(nc_out_rx_fast_clknb_aib1), .jtag_clkdr_in(clkdr_xr2l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_outpdir0_1),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_directinclkn[1]), .oclkn(oclkn_clkn1),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpoutp16 ( .idata1_in1_jtag_out(idat1_poutp16),
     .async_dat_in1_jtag_out(nc_async_dat_poutp16),
     .idata0_in1_jtag_out(idat0_poutp16),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp16),
     .prev_io_shift_en(rshift_en_poutp[14]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_pout[16]), .oclk_out(nc_oclk[16]),
     .oclkb_out(nc_oclkb[16]), .odat0_out(nc_odat0[16]),
     .odat1_out(nc_odat1[16]), .odat_async_out(nc_odat_async[16]),
     .pd_data_out(nc_pd_data[16]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp16),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[16]),
     .idata0_in1(idat0_poutp14), .idata1_in0(idat1[16]),
     .idata1_in1(idat1_poutp14), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[0]), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk_l[1]),
     .ilaunch_clk_in1(tx_launch_clk_l[1]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp16), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[16]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[16]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_poutp16),
     .odat1_aib(nc_odat1_aib_pout[16]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp16),
     .odat0_aib(nc_odat0_aib_pout[16]),
     .oclk_aib(nc_oclk_aib_pout[16]),
     .last_bs_out(nc_last_bs_out_poutp16),
     .oclkb_aib(nc_oclkb_aib_pout[16]), .jtag_clkdr_in(clkdr_xr5l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp14),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[16]), .oclkn(nc_oclkn_pout[16]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpoutp19 ( .idata1_in1_jtag_out(idat1_poutp19),
     .async_dat_in1_jtag_out(nc_async_dat_poutp19),
     .idata0_in1_jtag_out(idat0_poutp19),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp19),
     .prev_io_shift_en(rshift_en_poutp[17]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .dig_rstb(poutp_dig_rstb), .pd_data_aib(nc_pd_data_aib_pout[19]),
     .oclk_out(nc_oclk[19]), .oclkb_out(nc_oclkb[19]),
     .odat0_out(nc_odat0[19]), .odat1_out(nc_odat1[19]),
     .odat_async_out(nc_odat_async[19]), .pd_data_out(nc_pd_data[19]),
     .async_dat_in0(vssl_aibnd), .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp19),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[19]),
     .idata0_in1(idat0_poutp17), .idata1_in0(idat1[19]),
     .idata1_in1(idat1_poutp17), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[0]), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk_l[4]),
     .ilaunch_clk_in1(tx_launch_clk_l[4]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp19), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[19]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[19]), .pd_data_in1(vssl_aibnd),
     .jtag_clkdr_out(jtag_clkdr_out_poutp19),
     .odat1_aib(nc_odat1_aib_pout[19]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp19),
     .odat0_aib(nc_odat0_aib_pout[19]),
     .oclk_aib(nc_oclk_aib_pout[19]),
     .last_bs_out(nc_last_bs_out_poutp19),
     .oclkb_aib(nc_oclkb_aib_pout[19]), .jtag_clkdr_in(clkdr_xr6l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp17),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[19]), .oclkn(nc_oclkn_pout[19]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xasyncrx2 ( .idata1_in1_jtag_out(nc_idat1_async_in2),
     .async_dat_in1_jtag_out(nc_async_dat_async_in2),
     .idata0_in1_jtag_out(nc_idat0_async_in2),
     .jtag_clkdr_outn(jtag_clkdr_outn_inpshared2),
     .prev_io_shift_en(shift_en_ssrdout), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(output_rstb), .pd_data_aib(ncrx_pd_data_aib[2]),
     .oclk_out(odat_async[2]), .oclkb_out(ncrx_oclkb[2]),
     .odat0_out(ncrx_odat0[2]), .odat1_out(ncrx_odat1[2]),
     .odat_async_out(ncrx_async_data_out2),
     .pd_data_out(ncrx_pd_data[2]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(vssl_aibnd),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(idata0_ssrdout), .idata1_in0(vssl_aibnd),
     .idata1_in1(idata1_ssrdout), .idataselb_in0(vssl_aibnd),
     .idataselb_in1(idataselb_ssrdout), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(ilaunch_clk_ssrdout), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1(indrv_r34[1:0]), .ipdrv_in0({vssl_aibnd, vssl_aibnd}),
     .ipdrv_in1(ipdrv_r34[1:0]), .irxen_in0(irxen_r0[2:0]),
     .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(vssl_aibnd), .itxen_in1(itxen_ssrdout),
     .oclk_in1(oclk_inpshared0),
     .odat_async_aib(ncrx_odat_async_aib[2]),
     .oclkb_in1(oclkb_inpshared0), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_tx[2]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(avmm_sync_rstb), .jtag_clkdr_out(jtag_clkdr_async_in2),
     .odat1_aib(ncrx_odat1_aib[2]),
     .jtag_rx_scan_out(jtag_rx_scan_async_in2),
     .odat0_aib(ncrx_odat0_aib[2]), .oclk_aib(ncrx_oclk_aib2),
     .last_bs_out(nc_last_bs_out_diro2), .oclkb_aib(ncrx_oclkb_aib2),
     .jtag_clkdr_in(clkdr_xr3r), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_in_ssrdout),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_async_in[2]), .oclkn(ncrx_oclkn2),
     .iclkn(oclkn_inpshared3), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdirect_out2 (
     .idata1_in1_jtag_out(nc_idat1_outpdir3_1),
     .async_dat_in1_jtag_out(async_dat_outpdir3_1),
     .idata0_in1_jtag_out(nc_idat0_outpdir3_1),
     .jtag_clkdr_outn(jtag_clkdr_outn_outpdir3_1),
     .prev_io_shift_en(shift_en_in_chain2),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(ncdtx_pd_data_aib[2]), .oclk_out(ncdtx_oclk[2]),
     .oclkb_out(ncdtx_oclkb[2]), .odat0_out(ncdtx_odat0[2]),
     .odat1_out(ncdtx_odat1[2]), .odat_async_out(ncdtx_odat_async[2]),
     .pd_data_out(ncdtx_pd_data[2]),
     .async_dat_in0(idirectout_data[2]), .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(vssl_aibnd), .iclkin_dist_in1(vssl_aibnd),
     .idata0_in0(vssl_aibnd), .idata0_in1(vssl_aibnd),
     .idata1_in0(vssl_aibnd), .idata1_in1(vssl_aibnd),
     .idataselb_in0(idataselb[3]), .idataselb_in1(vssl_aibnd),
     .iddren_in0(vssl_aibnd), .iddren_in1(vssl_aibnd),
     .ilaunch_clk_in0(vssl_aibnd), .ilaunch_clk_in1(vssl_aibnd),
     .ilpbk_dat_in0(vssl_aibnd), .ilpbk_dat_in1(vssl_aibnd),
     .ilpbk_en_in0(vssl_aibnd), .ilpbk_en_in1(vssl_aibnd),
     .indrv_in0(indrv_r12[1:0]), .indrv_in1({vssl_aibnd, vssl_aibnd}),
     .ipdrv_in0(ipdrv_r12[1:0]), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .irxen_in1(irxen_in_chain2[2:0]), .istrbclk_in0(vssl_aibnd),
     .istrbclk_in1(vssl_aibnd), .itxen_in0(itxen[3]),
     .itxen_in1(vssl_aibnd), .oclk_in1(vssl_aibnd),
     .odat_async_aib(odirectin_data_out0_chain2),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_dtx[2]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(output_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_outpdir3_1),
     .odat1_aib(ncdtx_odat1_aib[2]),
     .jtag_rx_scan_out(jtag_rx_scan_out_outpdir3_1),
     .odat0_aib(ncdtx_odat0_aib[2]), .oclk_aib(oclk_outdir3_1),
     .last_bs_out(nc_last_bs_out_outpdir3_1),
     .oclkb_aib(oclkb_outdir3_1), .jtag_clkdr_in(clkdr_xr1r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_scan_in_chain2),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_directout[2]), .oclkn(ncdtx_oclkn[2]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpoutp17 ( .idata1_in1_jtag_out(idat1_poutp17),
     .async_dat_in1_jtag_out(nc_async_dat_poutp17),
     .idata0_in1_jtag_out(idat0_poutp17),
     .jtag_clkdr_outn(jtag_clkdr_outn_poutp17),
     .prev_io_shift_en(rshift_en_poutp[15]),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(nc_pd_data_aib_pout[17]), .oclk_out(nc_oclk[17]),
     .oclkb_out(nc_oclkb[17]), .odat0_out(nc_odat0[17]),
     .odat1_out(nc_odat1[17]), .odat_async_out(nc_odat_async[17]),
     .pd_data_out(nc_pd_data[17]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_poutp17),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0[17]),
     .idata0_in1(idat0_poutp15), .idata1_in0(idat1[17]),
     .idata1_in1(idat1_poutp15), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb[0]), .iddren_in0(iddren),
     .iddren_in1(iddren), .ilaunch_clk_in0(tx_launch_clk_l[0]),
     .ilaunch_clk_in1(tx_launch_clk_l[0]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_poutp17), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_aib_pout[17]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_poutp[17]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_poutp17),
     .odat1_aib(nc_odat1_aib_pout[17]),
     .jtag_rx_scan_out(jtag_rx_scan_out_poutp17),
     .odat0_aib(nc_odat0_aib_pout[17]),
     .oclk_aib(nc_oclk_aib_pout[17]),
     .last_bs_out(nc_last_bs_out_poutp17),
     .oclkb_aib(nc_oclkb_aib_pout[17]), .jtag_clkdr_in(clkdr_xr6l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_poutp15),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_dat[17]), .oclkn(nc_oclkn_pout[17]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xasynctx0 ( .idata1_in1_jtag_out(nc_idat1_async_out0),
     .async_dat_in1_jtag_out(async_dat_async_out0),
     .idata0_in1_jtag_out(nc_idat0_async_out0),
     .jtag_clkdr_outn(jtag_clkdr_outn_async_out0),
     .prev_io_shift_en(rshift_en_dtx[2]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(output_rstb), .pd_data_aib(nctx_pd_data_aib[0]),
     .oclk_out(nctx_oclk[0]), .oclkb_out(nctx_oclkb[0]),
     .odat0_out(nctx_odat0[0]), .odat1_out(nctx_odat1[0]),
     .odat_async_out(nctx_odat_async[0]),
     .pd_data_out(nctx_pd_data[0]), .async_dat_in0(iasyncdata[0]),
     .async_dat_in1(async_dat_outpdir3_1),
     .iclkin_dist_in0(vssl_aibnd), .iclkin_dist_in1(vssl_aibnd),
     .idata0_in0(vssl_aibnd), .idata0_in1(vssl_aibnd),
     .idata1_in0(vssl_aibnd), .idata1_in1(vssl_aibnd),
     .idataselb_in0(idataselb[2]), .idataselb_in1(idataselb[3]),
     .iddren_in0(vssl_aibnd), .iddren_in1(vssl_aibnd),
     .ilaunch_clk_in0(vssl_aibnd), .ilaunch_clk_in1(vssl_aibnd),
     .ilpbk_dat_in0(vssl_aibnd), .ilpbk_dat_in1(vssl_aibnd),
     .ilpbk_en_in0(vssl_aibnd), .ilpbk_en_in1(vssl_aibnd),
     .indrv_in0(indrv_r12[1:0]), .indrv_in1(indrv_r12[1:0]),
     .ipdrv_in0(ipdrv_r12[1:0]), .ipdrv_in1(ipdrv_r12[1:0]),
     .irxen_in0({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[2]), .itxen_in1(itxen[3]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(odat_async_oshared0), .oclkb_in1(vssl_aibnd),
     .odat0_in1(vssl_aibnd), .odat1_in1(vssl_aibnd),
     .odat_async_in1(odat_async_aib4), .shift_en(rshift_en_rx[0]),
     .pd_data_in1(vssl_aibnd), .dig_rstb(output_rstb),
     .jtag_clkdr_out(jtag_clkdr_async_out0),
     .odat1_aib(nctx_odat1_aib[0]),
     .jtag_rx_scan_out(jtag_rx_scan_async_out0),
     .odat0_aib(nctx_odat0_aib[0]), .oclk_aib(nctx_oclk_aib[0]),
     .last_bs_out(nc_last_bs_out_oshared0),
     .oclkb_aib(nctx_oclkb_aib[0]), .jtag_clkdr_in(clkdr_xr1r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_outpdir3_1),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_async_out[0]), .oclkn(nctx_oclkn[0]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdirect_out0 (
     .idata1_in1_jtag_out(nc_idat1_outpdir6),
     .async_dat_in1_jtag_out(idat0_outpdir6),
     .idata0_in1_jtag_out(nc_idat0_outpdir6),
     .jtag_clkdr_outn(jtag_clkdr_outn_outpdir6),
     .prev_io_shift_en(rshift_en_poutp[19]), .anlg_rstb(output_rstb),
     .pd_data_aib(ncdtx_pd_data_aib[0]), .oclk_out(ncdtx_oclk[0]),
     .oclkb_out(ncdtx_oclkb[0]), .odat0_out(ncdtx_odat0[0]),
     .odat1_out(ncdtx_odat1[0]), .odat_async_out(ncdtx_odat_async[0]),
     .pd_data_out(ncdtx_pd_data[0]),
     .async_dat_in0(idirectout_data[0]), .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(vssl_aibnd), .iclkin_dist_in1(vssl_aibnd),
     .idata0_in0(vssl_aibnd), .idata0_in1(idat0_poutp19),
     .idata1_in0(vssl_aibnd), .idata1_in1(idat1_poutp19),
     .idataselb_in0(idataselb[3]), .idataselb_in1(idataselb[0]),
     .iddren_in0(vssl_aibnd), .iddren_in1(iddren),
     .ilaunch_clk_in0(tx_launch_clk_l[8]),
     .ilaunch_clk_in1(tx_launch_clk_l[8]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[3]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(ncdtx_odat_async_aib[0]), .oclkb_in1(vssl_aibnd),
     .jtag_clksel(jtag_clksel), .odat0_in1(vssl_aibnd),
     .vssl_aibnd(vssl_aibnd), .odat1_in1(vssl_aibnd),
     .odat_async_in1(vssl_aibnd), .shift_en(rshift_en_dtx[0]),
     .pd_data_in1(vssl_aibnd), .dig_rstb(poutp_dig_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_outpdir6),
     .jtag_intest(jtag_intest), .odat1_aib(ncdtx_odat1_aib[0]),
     .jtag_rx_scan_out(jtag_rx_scan_out_outpdir6),
     .odat0_aib(ncdtx_odat0_aib[0]), .oclk_aib(ncdtx_oclk_aib0),
     .last_bs_out(nc_last_bs_out_outpdir6), .vccl_aibnd(vccl_aibnd),
     .oclkb_aib(ncdtx_oclkb_aib0), .jtag_clkdr_in(clkdr_xr6l),
     .jtag_rstb_en(jtag_rstb_en), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_poutp19),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_directout[0]), .oclkn(ncdtx_oclkn0),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdiin_clkp ( .idata1_in1_jtag_out(nc_idat1_dirclkp1),
     .async_dat_in1_jtag_out(nc_async_dat_dirclkp1),
     .idata0_in1_jtag_out(nc_idat0_dirclkp1),
     .jtag_clkdr_outn(jtag_clkdr_outn_inpclk0),
     .prev_io_shift_en(shift_en_outpclk1_1),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(output_rstb),
     .pd_data_aib(ncrx_pd_data_aib_clkp1),
     .oclk_out(out_rx_fast_clk[1]), .oclkb_out(out_rx_fast_clkb[1]),
     .odat0_out(nc_rxodat0_clkp[1]), .odat1_out(nc_rxodat1_clkp[1]),
     .odat_async_out(nc_rxodat_async_clkp[1]),
     .pd_data_out(nc_rxpd_data_clkp[1]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(async_dat_outpclk1_1),
     .iclkin_dist_in0(vssl_aibnd), .iclkin_dist_in1(vssl_aibnd),
     .idata0_in0(vssl_aibnd), .idata0_in1(vssl_aibnd),
     .idata1_in0(vssl_aibnd), .idata1_in1(vssl_aibnd),
     .idataselb_in0(vssl_aibnd), .idataselb_in1(idataselb_outpclk1_1),
     .iddren_in0(vssl_aibnd), .iddren_in1(vssl_aibnd),
     .ilaunch_clk_in0(vssl_aibnd), .ilaunch_clk_in1(vssl_aibnd),
     .ilpbk_dat_in0(vssl_aibnd), .ilpbk_dat_in1(vssl_aibnd),
     .ilpbk_en_in0(vssl_aibnd), .ilpbk_en_in1(vssl_aibnd),
     .indrv_in0({vssl_aibnd, vssl_aibnd}), .indrv_in1(indrv_r12[1:0]),
     .ipdrv_in0({vssl_aibnd, vssl_aibnd}), .ipdrv_in1(ipdrv_r12[1:0]),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .istrbclk_in0(vssl_aibnd),
     .istrbclk_in1(vssl_aibnd), .itxen_in0(vssl_aibnd),
     .itxen_in1(itxen_outpclk1_1), .oclk_in1(drx_oclk_aib[0]),
     .odat_async_aib(ncrx_odat_async_aib_clkp1),
     .oclkb_in1(drx_oclkb_aib[0]), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_dirclkp[1]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(output_rstb), .jtag_clkdr_out(jtag_clkdr_out_dirclkp1),
     .odat1_aib(nc_odat1_aib1),
     .jtag_rx_scan_out(jtag_rx_scan_out_dirclkp1),
     .odat0_aib(nc_odat0_aib1), .oclk_aib(nc_out_rx_fast_clk_aib1),
     .last_bs_out(nc_last_bs_out_inpclk0),
     .oclkb_aib(nc_out_rx_fast_clkb_aib1), .jtag_clkdr_in(clkdr_xr1l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_outpclk1_1),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_directinclkp[1]), .oclkn(nc_rxoclk_clkp1),
     .iclkn(oclkn_clkn1), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdirect_in1 ( .idata1_in1_jtag_out(nc_idat1_inpdir0),
     .async_dat_in1_jtag_out(nc_async_dat_inpdir0),
     .idata0_in1_jtag_out(nc_idat0_inpdir0),
     .jtag_clkdr_outn(jtag_clkdr_outn_inpdir0),
     .prev_io_shift_en(shift_en_pinp0), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(output_rstb), .pd_data_aib(ncdrx_pd_data_aib[1]),
     .oclk_out(ncdrx_oclk[1]), .oclkb_out(ncdrx_oclkb[1]),
     .odat0_out(ncdrx_odat0[1]), .odat1_out(ncdrx_odat1[1]),
     .odat_async_out(odirectin_data[1]),
     .pd_data_out(ncdrx_pd_data[1]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(iclkin_dist_pinp0),
     .iclkin_dist_in1(iclkin_dist_pinp0), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vssl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r1[2:0]), .irxen_in1(irxen_pinp0[2:0]),
     .istrbclk_in0(istrbclk_pinp0), .istrbclk_in1(istrbclk_pinp0),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(ncdrx_odat_async_aib[1]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(odat_async_chain2),
     .shift_en(rshift_en_drx[1]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(output_rstb), .jtag_clkdr_out(jtag_clkdr_out_chain2),
     .odat1_aib(odat1_inpdir0),
     .jtag_rx_scan_out(jtag_scan_out_chain2),
     .odat0_aib(odat0_inpdir0), .oclk_aib(ncdrx_oclk_aib[1]),
     .last_bs_out(nc_last_bs_out_inpdir0),
     .oclkb_aib(ncdrx_oclkb_aib[1]), .jtag_clkdr_in(clkdr_xr7r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_scan_pinp0),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_direct_input[1]), .oclkn(ncdrx_oclkn1),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top x750 ( .idata1_in1_jtag_out(nc_idat1_ptxclkin),
     .async_dat_in1_jtag_out(nc_async_dat_ptxclkin),
     .idata0_in1_jtag_out(nc_idat0_ptxclkin),
     .jtag_clkdr_outn(jtag_clkdr_outn_ptxclkin),
     .prev_io_shift_en(shift_en_voutp00), .anlg_rstb(output_rstb),
     .pd_data_aib(ncrx_pd_data_aib_clkp0),
     .oclk_out(nc_out_rx_fast_clk0_io), .oclkb_out(out_rx_fast_clkb[0]),
     .odat0_out(nc_rxodat0_clkp[0]), .odat1_out(nc_rxodat1_clkp[0]),
     .odat_async_out(nc_rxodat_async_clkp[0]),
     .pd_data_out(nc_rxpd_data_clkp[0]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(vssl_aibnd),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(idat0_voutp00), .idata1_in0(vssl_aibnd),
     .idata1_in1(idat1_voutp00), .idataselb_in0(vssl_aibnd),
     .idataselb_in1(idataselb_voutp00), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(ilaunch_clk_voutp00), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1(indrv_r34[1:0]), .ipdrv_in0({vssl_aibnd, vssl_aibnd}),
     .ipdrv_in1(ipdrv_r34[1:0]), .irxen_in0(irxen_r0[2:0]),
     .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(vssl_aibnd), .itxen_in1(itxen_voutp00),
     .oclk_in1(out_rx_fast_clk0_buf),
     .odat_async_aib(ncrx_odat_async_aib_clkp0),
     .oclkb_in1(oclkb_srclkout), .jtag_clksel(jtag_clksel),
     .odat0_in1(vssl_aibnd), .vssl_aibnd(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rshift_en_dirclkp[0]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(avmm_sync_rstb), .jtag_clkdr_out(jtag_clkdr_ptxclkin),
     .jtag_intest(jtag_intest), .odat1_aib(odat1_ptxclkin),
     .jtag_rx_scan_out(jtag_rx_scan_ptxclkin),
     .odat0_aib(odat0_ptxclkin), .oclk_aib(oclk_aib_ptxclkin),
     .last_bs_out(nc_last_bs_out_ptxclkin), .vccl_aibnd(vccl_aibnd),
     .oclkb_aib(oclkb_aib_ptxclkin), .jtag_clkdr_in(clkdr_xr3l),
     .jtag_rstb_en(jtag_rstb_en), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_voutp00),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_directinclkp[0]), .oclkn(nc_rxoclk_clkp0),
     .iclkn(oclkn_clkn0), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
assign outbuf_clk_buf = output_buffer_clk;

wire rb_dcc_byp_inv;
assign rb_dcc_byp_inv = ~rb_dcc_byp_dprio;

wire rb_dcc_en_dprio_buf , rb_dcc_manual_mode_dprio_buf;
assign rb_dcc_en_dprio_buf = rb_dcc_en_dprio;
assign rb_dcc_manual_mode_dprio_buf = rb_dcc_manual_mode_dprio ; //modified by Ana to pass linting(undriven),suspected typo[Nov4,2015]

aibnd_dcc_top  x711 ( .vcc_aibnd(vccl_aibnd),
     .rb_cont_cal(rb_dcc_manual_mode_dprio_buf), .scan_shift_n(scan_shift_n),
     .vss_aibnd(vssl_aibnd), .rb_clkdiv(rb_clkdiv[2:0]),
     .rb_dcc_manual_up(rb_dcc_manual_up[4:0]), .scan_rst_n(scan_rst_n),
     .clktree_out(clk_mimic0_buf),
     .rb_dcc_manual_dn(rb_dcc_manual_dn[4:0]),
     .dcc_dft_nrst_coding(dcc_dft_nrst_coding),
     .dcc_dft_nrst(dcc_dft_nrst), .dcc_dft_up(dcc_dft_up),
     .rb_dcc_dft(rb_dcc_dft), .rb_dcc_dft_sel(rb_dcc_dft_sel),
     .scan_out(dcc_scan_out), .scan_mode_n(scan_mode_n),
     .scan_in(scan_in), .pipeline_global_en(pipeline_global_en),
     .scan_clk_in(scan_clk_in), .rb_dcc_byp(rb_dcc_byp_inv),
     .vcc_io(vccl_aibnd), .clk_dcc(clktree_in), .dcc_done(dcc_done),
     .odll_dll2core(odcc_dll2core[12:0]), .clk_dcd(outbuf_clk_buf),
     .csr_reg(csr_reg[51:0]), .dcc_req(dcc_req),
     .idll_core2dll(oaibdftcore2dcc[2:0]), .idll_entest(idll_entest),
     .nfrzdrv(output_rstb), .rb_dcc_en(rb_dcc_en_dprio_buf),
     .rb_half_code(rb_half_code), .rb_selflock(rb_selflock),
     .test_clk_pll_en_n(rb_dcc_test_clk_pll_en_n));
aibnd_aliasd  aliasv8 ( .MINUS(ilaunch_clk_poutp18),      .PLUS(tx_launch_clk_l[9]));
aibnd_aliasd  aliasd21 ( .MINUS(shift_en_ptxclkinn),      .PLUS(rshift_en_dirclkn[0]));
aibnd_aliasd  aliasd20 ( .MINUS(oclkn_outpdir4_1), .PLUS(dtx_oclkn1));
aibnd_aliasd  aliasd12 ( .MINUS(shift_en_inpshared4),      .PLUS(rshift_en_rx[2]));
aibnd_aliasd  aliasd13 ( .MINUS(shift_en_oshared2), .PLUS(rshift_en_rx[3]));
aibnd_aliasd  aliasd18 ( .MINUS(shift_en_outpdir6), .PLUS(rshift_en_dtx[0]));
aibnd_aliasd  aliasv25[2:0] ( .MINUS(irxen_chain2[2:0]),      .PLUS(irxen_r1[2:0]));
aibnd_aliasd  aliasv24[2:0] ( .MINUS(irxen_inpdir3[2:0]),      .PLUS(irxen_r1[2:0]));
aibnd_aliasd  aliasv23[2:0] ( .MINUS(irxen_ptxclkin[2:0]),      .PLUS(irxen_r0[2:0]));
aibnd_aliasd  aliasd19 ( .MINUS(shift_en_poutp18),      .PLUS(rshift_en_poutp[18]));
aibnd_aliasd  aliasd17 ( .MINUS(shift_en_ptxclkin),      .PLUS(rshift_en_dirclkp[0]));
aibnd_aliasd  aliasd16 ( .MINUS(shift_en_outpdir1_1),      .PLUS(rshift_en_dtx[3]));
aibnd_aliasd  aliasd6 ( .MINUS(idataselb_oshared2), .PLUS(idataselb[2]));
aibnd_aliasd  aliasd9 ( .MINUS(itxen_oshared2), .PLUS(itxen[2]));
aibnd_aliasd  aliasd10[2:0] ( .MINUS(irxen_inpshared0[2:0]),      .PLUS(irxen_r0[2:0]));
aibnd_aliasd  aliasd3[2:0] ( .MINUS(irxen_inpshared4[2:0]),      .PLUS(irxen_r2[2:0]));
aibnd_aliasd  aliasv19[2:0] ( .MINUS(irxen_inpclk3[2:0]),      .PLUS(irxen_r1[2:0]));
aibnd_aliasd  aliasv15 ( .MINUS(idataselb_outpdir1_1), .PLUS(idataselb[3]));
aibnd_aliasd  aliasd11 ( .MINUS(shift_en_inpshared0),      .PLUS(rshift_en_tx[0]));
aibnd_aliasd  aliasd15 ( .MINUS(shift_en_inpclk0n),      .PLUS(rshift_en_dirclkn[1]));
aibnd_aliasd  aliasv12 ( .MINUS(itxen_outpdir1_1), .PLUS(itxen[3]));
aibnd_aliasd  aliasv7 ( .MINUS(itxen_outpdir6), .PLUS(itxen[3]));
aibnd_aliasd  aliasv9 ( .MINUS(idataselb_poutp18), .PLUS(idataselb[0]));
aibnd_aliasd  aliasv17 ( .MINUS(iddren_poutp18), .PLUS(iddren));
aibnd_aliasd  aliasd23 ( .MINUS(shift_en_inpclk3), .PLUS(rshift_en_drx[2]));
aibnd_aliasd  aliasd22 ( .MINUS(shift_en_out_chain2),      .PLUS(rshift_en_drx[1]));
aibnd_aliasd  aliasv16 ( .MINUS(idataselb_outpdir6), .PLUS(idataselb[3]));
aibnd_aliasd  aliasv1 ( .MINUS(itxen_poutp18), .PLUS(itxen[0]));
aibnd_aliasd  aliasd14 ( .MINUS(shift_en_inpdir3), .PLUS(rshift_en_drx[0]));

aibnd_clkmux2 xtx_rx_clkmx ( 
      .oclk_out(out_rx_fast_clk[0]),
     .mux_sel(rshift_en_dirclkp[0]), .oclk_in0(oclk_aib_ptxclkin),
     .oclk_in1(oclk_srclkout));

assign out_rx_fast_clk0_buf = out_rx_fast_clk[0] ;

assign oaibdftdll2core[10] = mux_dft_dll2core[10];
assign oaibdftdll2core[11] = mux_dft_dll2core[11];
assign oaibdftdll2core[9] = mux_dft_dll2core[9];
assign buf_dcc2core[1] = odcc_dll2core[1];
assign oaibdftdll2core[12] = mux_dft_dll2core[12];
assign oaibdftcore2dll[2] = oaibdftcore2dcc[2];
assign oaibdftcore2dcc[1] = iaibdftcore2dll[1];
assign buf_dcc2core[2] = odcc_dll2core[2];
assign oaibdftcore2dll[1] = oaibdftcore2dcc[1];
assign buf_dcc2core[11] = odcc_dll2core[11];
assign buf_dll2core[8] = idll_dll2core[8];
assign buf_dll2core[7] = idll_dll2core[7];
assign buf_dll2core[5] = idll_dll2core[5];
assign oaibdftdll2core[8] = mux_dft_dll2core[8];
assign buf_dcc2core[6] = odcc_dll2core[6];
assign oaibdftdll2core[7] = mux_dft_dll2core[7];
assign buf_dcc2core[8] = odcc_dll2core[8];
assign buf_dll2core[6] = idll_dll2core[6];
assign oaibdftdll2core[5] = mux_dft_dll2core[5];
assign buf_dcc2core[7] = odcc_dll2core[7];
assign oaibdftdll2core[6] = mux_dft_dll2core[6];
assign buf_dcc2core[5] = odcc_dll2core[5];
assign buf_dll2core[4] = idll_dll2core[4];
assign buf_dcc2core[12] = odcc_dll2core[12];
assign buf_dll2core[10] = idll_dll2core[10];
assign buf_dll2core[9] = idll_dll2core[9];
assign buf_dll2core[11] = idll_dll2core[11];
assign oaibdftdll2core[4] = mux_dft_dll2core[4];
assign buf_dcc2core[4] = odcc_dll2core[4];
assign buf_dcc2core[3] = odcc_dll2core[3];
assign oaibdftdll2core[0] = mux_dft_dll2core[0];
assign buf_dcc2core[0] = odcc_dll2core[0];
assign oaibdftcore2dcc[2] = iaibdftcore2dll[2];
assign buf_dll2core[1] = idll_dll2core[1];
assign oaibdftdll2core[1] = mux_dft_dll2core[1];
assign oaibdftcore2dll[0] = oaibdftcore2dcc[0];
assign buf_dll2core[0] = idll_dll2core[0];
assign oaibdftcore2dcc[0] = iaibdftcore2dll[0];
assign buf_dcc2core[9] = odcc_dll2core[9];
assign buf_dll2core[12] = idll_dll2core[12];
assign oaibdftdll2core[2] = mux_dft_dll2core[2];
assign buf_dll2core[2] = idll_dll2core[2];
assign buf_dll2core[3] = idll_dll2core[3];
assign oaibdftdll2core[3] = mux_dft_dll2core[3];
assign buf_dcc2core[10] = odcc_dll2core[10];
assign mux_dft_dll2core[2] = rb_dcc_dll_dft_sel ? buf_dcc2core[2] : buf_dll2core[2];
assign mux_dft_dll2core[10] = rb_dcc_dll_dft_sel ? buf_dcc2core[10] : buf_dll2core[10];
assign mux_dft_dll2core[6] = rb_dcc_dll_dft_sel ? buf_dcc2core[6] : buf_dll2core[6];
assign mux_dft_dll2core[8] = rb_dcc_dll_dft_sel ? buf_dcc2core[8] : buf_dll2core[8];
assign mux_dft_dll2core[7] = rb_dcc_dll_dft_sel ? buf_dcc2core[7] : buf_dll2core[7];
assign mux_dft_dll2core[5] = rb_dcc_dll_dft_sel ? buf_dcc2core[5] : buf_dll2core[5];
assign mux_dft_dll2core[4] = rb_dcc_dll_dft_sel ? buf_dcc2core[4] : buf_dll2core[4];
assign mux_dft_dll2core[3] = rb_dcc_dll_dft_sel ? buf_dcc2core[3] : buf_dll2core[3];
assign mux_dft_dll2core[0] = rb_dcc_dll_dft_sel ? buf_dcc2core[0] : buf_dll2core[0];
assign mux_dft_dll2core[1] = rb_dcc_dll_dft_sel ? buf_dcc2core[1] : buf_dll2core[1];
assign mux_dft_dll2core[9] = rb_dcc_dll_dft_sel ? buf_dcc2core[9] : buf_dll2core[9];
assign mux_dft_dll2core[12] = rb_dcc_dll_dft_sel ? buf_dcc2core[12] : buf_dll2core[12];
assign mux_dft_dll2core[11] = rb_dcc_dll_dft_sel ? buf_dcc2core[11] : buf_dll2core[11];
assign scan_out = dcc_scan_out;
//assign clk_mimic0_buf = clk_mimic0;
assign clk_mimic0_buf = 1'b0;
assign clk_mimic1_buf = clk_mimic1;
assign dft_rx_clk = gated_clk_mimic1;
assign gated_clk_mimic1 = clk_mimic1_buf & dll_csr_reg6;
assign nc_clk_repb = !clk_rep;
//assign nc_clk_mimic = !clk_mimic;
assign nc_clk_mimic = 1'b1;


endmodule

