// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. 
//------------------------------------------------------------------------
// Copyright (c) 2012 Altera Corporation. .
module aibndaux_aliasd ( PLUS, MINUS );

	input   PLUS;
	output  MINUS;

	assign MINUS = PLUS;

endmodule





