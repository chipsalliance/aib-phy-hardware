// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. All rights reserved
module aibnd_aliasv ( .PLUS(w), .MINUS(w) );

	inout   w;
	wire    w;

endmodule





