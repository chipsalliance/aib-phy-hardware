// =====================================================================================
//
// Description: Verilog Nestlist
//   Component: 16 channel EMIB between master AIB model and FPGA AIB slave
//        date: 10/28/2020
//
// =====================================================================================
 module emib (
// ## START OF  ch0 ( ##
        inout [95:0] m0_ch0_aib,
 	inout  nd_aib95_ch0_x0y0, 
	inout  nd_aib94_ch0_x0y0, 
	inout  nd_aib93_ch0_x0y0, 
	inout  nd_aib92_ch0_x0y0, 
	inout  nd_aib91_ch0_x0y0, 
	inout  nd_aib90_ch0_x0y0, 
	inout  nd_aib89_ch0_x0y0, 
	inout  nd_aib88_ch0_x0y0, 
	inout  nd_aib87_ch0_x0y0, 
	inout  nd_aib86_ch0_x0y0, 
	inout  nd_aib85_ch0_x0y0, 
	inout  nd_aib84_ch0_x0y0, 
	inout  nd_aib83_ch0_x0y0, 
	inout  nd_aib82_ch0_x0y0, 
	inout  nd_aib81_ch0_x0y0, 
	inout  nd_aib80_ch0_x0y0, 
	inout  nd_aib79_ch0_x0y0, 
	inout  nd_aib78_ch0_x0y0, 
	inout  nd_aib77_ch0_x0y0, 
	inout  nd_aib76_ch0_x0y0, 
	inout  nd_aib75_ch0_x0y0, 
	inout  nd_aib74_ch0_x0y0, 
	inout  nd_aib73_ch0_x0y0, 
	inout  nd_aib72_ch0_x0y0, 
	inout  nd_aib71_ch0_x0y0, 
	inout  nd_aib70_ch0_x0y0, 
	inout  nd_aib69_ch0_x0y0, 
	inout  nd_aib68_ch0_x0y0, 
	inout  nd_aib67_ch0_x0y0, 
	inout  nd_aib66_ch0_x0y0, 
	inout  nd_aib65_ch0_x0y0, 
	inout  nd_aib64_ch0_x0y0, 
	inout  nd_aib63_ch0_x0y0, 
	inout  nd_aib62_ch0_x0y0, 
	inout  nd_aib61_ch0_x0y0, 
	inout  nd_aib60_ch0_x0y0, 
	inout  nd_aib59_ch0_x0y0, 
	inout  nd_aib58_ch0_x0y0, 
	inout  nd_aib57_ch0_x0y0, 
	inout  nd_aib56_ch0_x0y0, 
	inout  nd_aib55_ch0_x0y0, 
	inout  nd_aib54_ch0_x0y0, 
	inout  nd_aib53_ch0_x0y0, 
	inout  nd_aib52_ch0_x0y0, 
	inout  nd_aib51_ch0_x0y0, 
	inout  nd_aib50_ch0_x0y0, 
	inout  nd_aib49_ch0_x0y0, 
	inout  nd_aib48_ch0_x0y0, 
	inout  nd_aib47_ch0_x0y0, 
	inout  nd_aib46_ch0_x0y0, 
	inout  nd_aib45_ch0_x0y0, 
	inout  nd_aib44_ch0_x0y0, 
	inout  nd_aib43_ch0_x0y0, 
	inout  nd_aib42_ch0_x0y0, 
	inout  nd_aib41_ch0_x0y0, 
	inout  nd_aib40_ch0_x0y0, 
	inout  nd_aib39_ch0_x0y0, 
	inout  nd_aib38_ch0_x0y0, 
	inout  nd_aib37_ch0_x0y0, 
	inout  nd_aib36_ch0_x0y0, 
	inout  nd_aib35_ch0_x0y0, 
	inout  nd_aib34_ch0_x0y0, 
	inout  nd_aib33_ch0_x0y0, 
	inout  nd_aib32_ch0_x0y0, 
	inout  nd_aib31_ch0_x0y0, 
	inout  nd_aib30_ch0_x0y0, 
	inout  nd_aib29_ch0_x0y0, 
	inout  nd_aib28_ch0_x0y0, 
	inout  nd_aib27_ch0_x0y0, 
	inout  nd_aib26_ch0_x0y0, 
	inout  nd_aib25_ch0_x0y0, 
	inout  nd_aib24_ch0_x0y0, 
	inout  nd_aib23_ch0_x0y0, 
	inout  nd_aib22_ch0_x0y0, 
	inout  nd_aib21_ch0_x0y0, 
	inout  nd_aib20_ch0_x0y0, 
	inout  nd_aib19_ch0_x0y0, 
	inout  nd_aib18_ch0_x0y0, 
	inout  nd_aib17_ch0_x0y0, 
	inout  nd_aib16_ch0_x0y0, 
	inout  nd_aib15_ch0_x0y0, 
	inout  nd_aib14_ch0_x0y0, 
	inout  nd_aib13_ch0_x0y0, 
	inout  nd_aib12_ch0_x0y0, 
	inout  nd_aib11_ch0_x0y0, 
	inout  nd_aib10_ch0_x0y0, 
	inout  nd_aib9_ch0_x0y0, 
	inout  nd_aib8_ch0_x0y0, 
	inout  nd_aib7_ch0_x0y0, 
	inout  nd_aib6_ch0_x0y0, 
	inout  nd_aib5_ch0_x0y0, 
	inout  nd_aib4_ch0_x0y0, 
	inout  nd_aib3_ch0_x0y0, 
	inout  nd_aib2_ch0_x0y0, 
	inout  nd_aib1_ch0_x0y0, 
	inout  nd_aib0_ch0_x0y0, 
// ## START OF  ch1 ( ##
        inout [95:0] m0_ch1_aib,
 	inout  nd_aib95_ch1_x0y0, 
	inout  nd_aib94_ch1_x0y0, 
	inout  nd_aib93_ch1_x0y0, 
	inout  nd_aib92_ch1_x0y0, 
	inout  nd_aib91_ch1_x0y0, 
	inout  nd_aib90_ch1_x0y0, 
	inout  nd_aib89_ch1_x0y0, 
	inout  nd_aib88_ch1_x0y0, 
	inout  nd_aib87_ch1_x0y0, 
	inout  nd_aib86_ch1_x0y0, 
	inout  nd_aib85_ch1_x0y0, 
	inout  nd_aib84_ch1_x0y0, 
	inout  nd_aib83_ch1_x0y0, 
	inout  nd_aib82_ch1_x0y0, 
	inout  nd_aib81_ch1_x0y0, 
	inout  nd_aib80_ch1_x0y0, 
	inout  nd_aib79_ch1_x0y0, 
	inout  nd_aib78_ch1_x0y0, 
	inout  nd_aib77_ch1_x0y0, 
	inout  nd_aib76_ch1_x0y0, 
	inout  nd_aib75_ch1_x0y0, 
	inout  nd_aib74_ch1_x0y0, 
	inout  nd_aib73_ch1_x0y0, 
	inout  nd_aib72_ch1_x0y0, 
	inout  nd_aib71_ch1_x0y0, 
	inout  nd_aib70_ch1_x0y0, 
	inout  nd_aib69_ch1_x0y0, 
	inout  nd_aib68_ch1_x0y0, 
	inout  nd_aib67_ch1_x0y0, 
	inout  nd_aib66_ch1_x0y0, 
	inout  nd_aib65_ch1_x0y0, 
	inout  nd_aib64_ch1_x0y0, 
	inout  nd_aib63_ch1_x0y0, 
	inout  nd_aib62_ch1_x0y0, 
	inout  nd_aib61_ch1_x0y0, 
	inout  nd_aib60_ch1_x0y0, 
	inout  nd_aib59_ch1_x0y0, 
	inout  nd_aib58_ch1_x0y0, 
	inout  nd_aib57_ch1_x0y0, 
	inout  nd_aib56_ch1_x0y0, 
	inout  nd_aib55_ch1_x0y0, 
	inout  nd_aib54_ch1_x0y0, 
	inout  nd_aib53_ch1_x0y0, 
	inout  nd_aib52_ch1_x0y0, 
	inout  nd_aib51_ch1_x0y0, 
	inout  nd_aib50_ch1_x0y0, 
	inout  nd_aib49_ch1_x0y0, 
	inout  nd_aib48_ch1_x0y0, 
	inout  nd_aib47_ch1_x0y0, 
	inout  nd_aib46_ch1_x0y0, 
	inout  nd_aib45_ch1_x0y0, 
	inout  nd_aib44_ch1_x0y0, 
	inout  nd_aib43_ch1_x0y0, 
	inout  nd_aib42_ch1_x0y0, 
	inout  nd_aib41_ch1_x0y0, 
	inout  nd_aib40_ch1_x0y0, 
	inout  nd_aib39_ch1_x0y0, 
	inout  nd_aib38_ch1_x0y0, 
	inout  nd_aib37_ch1_x0y0, 
	inout  nd_aib36_ch1_x0y0, 
	inout  nd_aib35_ch1_x0y0, 
	inout  nd_aib34_ch1_x0y0, 
	inout  nd_aib33_ch1_x0y0, 
	inout  nd_aib32_ch1_x0y0, 
	inout  nd_aib31_ch1_x0y0, 
	inout  nd_aib30_ch1_x0y0, 
	inout  nd_aib29_ch1_x0y0, 
	inout  nd_aib28_ch1_x0y0, 
	inout  nd_aib27_ch1_x0y0, 
	inout  nd_aib26_ch1_x0y0, 
	inout  nd_aib25_ch1_x0y0, 
	inout  nd_aib24_ch1_x0y0, 
	inout  nd_aib23_ch1_x0y0, 
	inout  nd_aib22_ch1_x0y0, 
	inout  nd_aib21_ch1_x0y0, 
	inout  nd_aib20_ch1_x0y0, 
	inout  nd_aib19_ch1_x0y0, 
	inout  nd_aib18_ch1_x0y0, 
	inout  nd_aib17_ch1_x0y0, 
	inout  nd_aib16_ch1_x0y0, 
	inout  nd_aib15_ch1_x0y0, 
	inout  nd_aib14_ch1_x0y0, 
	inout  nd_aib13_ch1_x0y0, 
	inout  nd_aib12_ch1_x0y0, 
	inout  nd_aib11_ch1_x0y0, 
	inout  nd_aib10_ch1_x0y0, 
	inout  nd_aib9_ch1_x0y0, 
	inout  nd_aib8_ch1_x0y0, 
	inout  nd_aib7_ch1_x0y0, 
	inout  nd_aib6_ch1_x0y0, 
	inout  nd_aib5_ch1_x0y0, 
	inout  nd_aib4_ch1_x0y0, 
	inout  nd_aib3_ch1_x0y0, 
	inout  nd_aib2_ch1_x0y0, 
	inout  nd_aib1_ch1_x0y0, 
	inout  nd_aib0_ch1_x0y0, 
// ## START OF  ch2 ( ##
        inout [95:0] m0_ch2_aib,
 	inout  nd_aib95_ch2_x0y0, 
	inout  nd_aib94_ch2_x0y0, 
	inout  nd_aib93_ch2_x0y0, 
	inout  nd_aib92_ch2_x0y0, 
	inout  nd_aib91_ch2_x0y0, 
	inout  nd_aib90_ch2_x0y0, 
	inout  nd_aib89_ch2_x0y0, 
	inout  nd_aib88_ch2_x0y0, 
	inout  nd_aib87_ch2_x0y0, 
	inout  nd_aib86_ch2_x0y0, 
	inout  nd_aib85_ch2_x0y0, 
	inout  nd_aib84_ch2_x0y0, 
	inout  nd_aib83_ch2_x0y0, 
	inout  nd_aib82_ch2_x0y0, 
	inout  nd_aib81_ch2_x0y0, 
	inout  nd_aib80_ch2_x0y0, 
	inout  nd_aib79_ch2_x0y0, 
	inout  nd_aib78_ch2_x0y0, 
	inout  nd_aib77_ch2_x0y0, 
	inout  nd_aib76_ch2_x0y0, 
	inout  nd_aib75_ch2_x0y0, 
	inout  nd_aib74_ch2_x0y0, 
	inout  nd_aib73_ch2_x0y0, 
	inout  nd_aib72_ch2_x0y0, 
	inout  nd_aib71_ch2_x0y0, 
	inout  nd_aib70_ch2_x0y0, 
	inout  nd_aib69_ch2_x0y0, 
	inout  nd_aib68_ch2_x0y0, 
	inout  nd_aib67_ch2_x0y0, 
	inout  nd_aib66_ch2_x0y0, 
	inout  nd_aib65_ch2_x0y0, 
	inout  nd_aib64_ch2_x0y0, 
	inout  nd_aib63_ch2_x0y0, 
	inout  nd_aib62_ch2_x0y0, 
	inout  nd_aib61_ch2_x0y0, 
	inout  nd_aib60_ch2_x0y0, 
	inout  nd_aib59_ch2_x0y0, 
	inout  nd_aib58_ch2_x0y0, 
	inout  nd_aib57_ch2_x0y0, 
	inout  nd_aib56_ch2_x0y0, 
	inout  nd_aib55_ch2_x0y0, 
	inout  nd_aib54_ch2_x0y0, 
	inout  nd_aib53_ch2_x0y0, 
	inout  nd_aib52_ch2_x0y0, 
	inout  nd_aib51_ch2_x0y0, 
	inout  nd_aib50_ch2_x0y0, 
	inout  nd_aib49_ch2_x0y0, 
	inout  nd_aib48_ch2_x0y0, 
	inout  nd_aib47_ch2_x0y0, 
	inout  nd_aib46_ch2_x0y0, 
	inout  nd_aib45_ch2_x0y0, 
	inout  nd_aib44_ch2_x0y0, 
	inout  nd_aib43_ch2_x0y0, 
	inout  nd_aib42_ch2_x0y0, 
	inout  nd_aib41_ch2_x0y0, 
	inout  nd_aib40_ch2_x0y0, 
	inout  nd_aib39_ch2_x0y0, 
	inout  nd_aib38_ch2_x0y0, 
	inout  nd_aib37_ch2_x0y0, 
	inout  nd_aib36_ch2_x0y0, 
	inout  nd_aib35_ch2_x0y0, 
	inout  nd_aib34_ch2_x0y0, 
	inout  nd_aib33_ch2_x0y0, 
	inout  nd_aib32_ch2_x0y0, 
	inout  nd_aib31_ch2_x0y0, 
	inout  nd_aib30_ch2_x0y0, 
	inout  nd_aib29_ch2_x0y0, 
	inout  nd_aib28_ch2_x0y0, 
	inout  nd_aib27_ch2_x0y0, 
	inout  nd_aib26_ch2_x0y0, 
	inout  nd_aib25_ch2_x0y0, 
	inout  nd_aib24_ch2_x0y0, 
	inout  nd_aib23_ch2_x0y0, 
	inout  nd_aib22_ch2_x0y0, 
	inout  nd_aib21_ch2_x0y0, 
	inout  nd_aib20_ch2_x0y0, 
	inout  nd_aib19_ch2_x0y0, 
	inout  nd_aib18_ch2_x0y0, 
	inout  nd_aib17_ch2_x0y0, 
	inout  nd_aib16_ch2_x0y0, 
	inout  nd_aib15_ch2_x0y0, 
	inout  nd_aib14_ch2_x0y0, 
	inout  nd_aib13_ch2_x0y0, 
	inout  nd_aib12_ch2_x0y0, 
	inout  nd_aib11_ch2_x0y0, 
	inout  nd_aib10_ch2_x0y0, 
	inout  nd_aib9_ch2_x0y0, 
	inout  nd_aib8_ch2_x0y0, 
	inout  nd_aib7_ch2_x0y0, 
	inout  nd_aib6_ch2_x0y0, 
	inout  nd_aib5_ch2_x0y0, 
	inout  nd_aib4_ch2_x0y0, 
	inout  nd_aib3_ch2_x0y0, 
	inout  nd_aib2_ch2_x0y0, 
	inout  nd_aib1_ch2_x0y0, 
	inout  nd_aib0_ch2_x0y0, 
// ## START OF  ch3 ( ##
        inout [95:0] m0_ch3_aib,
 	inout  nd_aib95_ch3_x0y0, 
	inout  nd_aib94_ch3_x0y0, 
	inout  nd_aib93_ch3_x0y0, 
	inout  nd_aib92_ch3_x0y0, 
	inout  nd_aib91_ch3_x0y0, 
	inout  nd_aib90_ch3_x0y0, 
	inout  nd_aib89_ch3_x0y0, 
	inout  nd_aib88_ch3_x0y0, 
	inout  nd_aib87_ch3_x0y0, 
	inout  nd_aib86_ch3_x0y0, 
	inout  nd_aib85_ch3_x0y0, 
	inout  nd_aib84_ch3_x0y0, 
	inout  nd_aib83_ch3_x0y0, 
	inout  nd_aib82_ch3_x0y0, 
	inout  nd_aib81_ch3_x0y0, 
	inout  nd_aib80_ch3_x0y0, 
	inout  nd_aib79_ch3_x0y0, 
	inout  nd_aib78_ch3_x0y0, 
	inout  nd_aib77_ch3_x0y0, 
	inout  nd_aib76_ch3_x0y0, 
	inout  nd_aib75_ch3_x0y0, 
	inout  nd_aib74_ch3_x0y0, 
	inout  nd_aib73_ch3_x0y0, 
	inout  nd_aib72_ch3_x0y0, 
	inout  nd_aib71_ch3_x0y0, 
	inout  nd_aib70_ch3_x0y0, 
	inout  nd_aib69_ch3_x0y0, 
	inout  nd_aib68_ch3_x0y0, 
	inout  nd_aib67_ch3_x0y0, 
	inout  nd_aib66_ch3_x0y0, 
	inout  nd_aib65_ch3_x0y0, 
	inout  nd_aib64_ch3_x0y0, 
	inout  nd_aib63_ch3_x0y0, 
	inout  nd_aib62_ch3_x0y0, 
	inout  nd_aib61_ch3_x0y0, 
	inout  nd_aib60_ch3_x0y0, 
	inout  nd_aib59_ch3_x0y0, 
	inout  nd_aib58_ch3_x0y0, 
	inout  nd_aib57_ch3_x0y0, 
	inout  nd_aib56_ch3_x0y0, 
	inout  nd_aib55_ch3_x0y0, 
	inout  nd_aib54_ch3_x0y0, 
	inout  nd_aib53_ch3_x0y0, 
	inout  nd_aib52_ch3_x0y0, 
	inout  nd_aib51_ch3_x0y0, 
	inout  nd_aib50_ch3_x0y0, 
	inout  nd_aib49_ch3_x0y0, 
	inout  nd_aib48_ch3_x0y0, 
	inout  nd_aib47_ch3_x0y0, 
	inout  nd_aib46_ch3_x0y0, 
	inout  nd_aib45_ch3_x0y0, 
	inout  nd_aib44_ch3_x0y0, 
	inout  nd_aib43_ch3_x0y0, 
	inout  nd_aib42_ch3_x0y0, 
	inout  nd_aib41_ch3_x0y0, 
	inout  nd_aib40_ch3_x0y0, 
	inout  nd_aib39_ch3_x0y0, 
	inout  nd_aib38_ch3_x0y0, 
	inout  nd_aib37_ch3_x0y0, 
	inout  nd_aib36_ch3_x0y0, 
	inout  nd_aib35_ch3_x0y0, 
	inout  nd_aib34_ch3_x0y0, 
	inout  nd_aib33_ch3_x0y0, 
	inout  nd_aib32_ch3_x0y0, 
	inout  nd_aib31_ch3_x0y0, 
	inout  nd_aib30_ch3_x0y0, 
	inout  nd_aib29_ch3_x0y0, 
	inout  nd_aib28_ch3_x0y0, 
	inout  nd_aib27_ch3_x0y0, 
	inout  nd_aib26_ch3_x0y0, 
	inout  nd_aib25_ch3_x0y0, 
	inout  nd_aib24_ch3_x0y0, 
	inout  nd_aib23_ch3_x0y0, 
	inout  nd_aib22_ch3_x0y0, 
	inout  nd_aib21_ch3_x0y0, 
	inout  nd_aib20_ch3_x0y0, 
	inout  nd_aib19_ch3_x0y0, 
	inout  nd_aib18_ch3_x0y0, 
	inout  nd_aib17_ch3_x0y0, 
	inout  nd_aib16_ch3_x0y0, 
	inout  nd_aib15_ch3_x0y0, 
	inout  nd_aib14_ch3_x0y0, 
	inout  nd_aib13_ch3_x0y0, 
	inout  nd_aib12_ch3_x0y0, 
	inout  nd_aib11_ch3_x0y0, 
	inout  nd_aib10_ch3_x0y0, 
	inout  nd_aib9_ch3_x0y0, 
	inout  nd_aib8_ch3_x0y0, 
	inout  nd_aib7_ch3_x0y0, 
	inout  nd_aib6_ch3_x0y0, 
	inout  nd_aib5_ch3_x0y0, 
	inout  nd_aib4_ch3_x0y0, 
	inout  nd_aib3_ch3_x0y0, 
	inout  nd_aib2_ch3_x0y0, 
	inout  nd_aib1_ch3_x0y0, 
	inout  nd_aib0_ch3_x0y0, 
// ## START OF  ch4 ( ##
        inout [95:0] m0_ch4_aib,
 	inout  nd_aib95_ch4_x0y0, 
	inout  nd_aib94_ch4_x0y0, 
	inout  nd_aib93_ch4_x0y0, 
	inout  nd_aib92_ch4_x0y0, 
	inout  nd_aib91_ch4_x0y0, 
	inout  nd_aib90_ch4_x0y0, 
	inout  nd_aib89_ch4_x0y0, 
	inout  nd_aib88_ch4_x0y0, 
	inout  nd_aib87_ch4_x0y0, 
	inout  nd_aib86_ch4_x0y0, 
	inout  nd_aib85_ch4_x0y0, 
	inout  nd_aib84_ch4_x0y0, 
	inout  nd_aib83_ch4_x0y0, 
	inout  nd_aib82_ch4_x0y0, 
	inout  nd_aib81_ch4_x0y0, 
	inout  nd_aib80_ch4_x0y0, 
	inout  nd_aib79_ch4_x0y0, 
	inout  nd_aib78_ch4_x0y0, 
	inout  nd_aib77_ch4_x0y0, 
	inout  nd_aib76_ch4_x0y0, 
	inout  nd_aib75_ch4_x0y0, 
	inout  nd_aib74_ch4_x0y0, 
	inout  nd_aib73_ch4_x0y0, 
	inout  nd_aib72_ch4_x0y0, 
	inout  nd_aib71_ch4_x0y0, 
	inout  nd_aib70_ch4_x0y0, 
	inout  nd_aib69_ch4_x0y0, 
	inout  nd_aib68_ch4_x0y0, 
	inout  nd_aib67_ch4_x0y0, 
	inout  nd_aib66_ch4_x0y0, 
	inout  nd_aib65_ch4_x0y0, 
	inout  nd_aib64_ch4_x0y0, 
	inout  nd_aib63_ch4_x0y0, 
	inout  nd_aib62_ch4_x0y0, 
	inout  nd_aib61_ch4_x0y0, 
	inout  nd_aib60_ch4_x0y0, 
	inout  nd_aib59_ch4_x0y0, 
	inout  nd_aib58_ch4_x0y0, 
	inout  nd_aib57_ch4_x0y0, 
	inout  nd_aib56_ch4_x0y0, 
	inout  nd_aib55_ch4_x0y0, 
	inout  nd_aib54_ch4_x0y0, 
	inout  nd_aib53_ch4_x0y0, 
	inout  nd_aib52_ch4_x0y0, 
	inout  nd_aib51_ch4_x0y0, 
	inout  nd_aib50_ch4_x0y0, 
	inout  nd_aib49_ch4_x0y0, 
	inout  nd_aib48_ch4_x0y0, 
	inout  nd_aib47_ch4_x0y0, 
	inout  nd_aib46_ch4_x0y0, 
	inout  nd_aib45_ch4_x0y0, 
	inout  nd_aib44_ch4_x0y0, 
	inout  nd_aib43_ch4_x0y0, 
	inout  nd_aib42_ch4_x0y0, 
	inout  nd_aib41_ch4_x0y0, 
	inout  nd_aib40_ch4_x0y0, 
	inout  nd_aib39_ch4_x0y0, 
	inout  nd_aib38_ch4_x0y0, 
	inout  nd_aib37_ch4_x0y0, 
	inout  nd_aib36_ch4_x0y0, 
	inout  nd_aib35_ch4_x0y0, 
	inout  nd_aib34_ch4_x0y0, 
	inout  nd_aib33_ch4_x0y0, 
	inout  nd_aib32_ch4_x0y0, 
	inout  nd_aib31_ch4_x0y0, 
	inout  nd_aib30_ch4_x0y0, 
	inout  nd_aib29_ch4_x0y0, 
	inout  nd_aib28_ch4_x0y0, 
	inout  nd_aib27_ch4_x0y0, 
	inout  nd_aib26_ch4_x0y0, 
	inout  nd_aib25_ch4_x0y0, 
	inout  nd_aib24_ch4_x0y0, 
	inout  nd_aib23_ch4_x0y0, 
	inout  nd_aib22_ch4_x0y0, 
	inout  nd_aib21_ch4_x0y0, 
	inout  nd_aib20_ch4_x0y0, 
	inout  nd_aib19_ch4_x0y0, 
	inout  nd_aib18_ch4_x0y0, 
	inout  nd_aib17_ch4_x0y0, 
	inout  nd_aib16_ch4_x0y0, 
	inout  nd_aib15_ch4_x0y0, 
	inout  nd_aib14_ch4_x0y0, 
	inout  nd_aib13_ch4_x0y0, 
	inout  nd_aib12_ch4_x0y0, 
	inout  nd_aib11_ch4_x0y0, 
	inout  nd_aib10_ch4_x0y0, 
	inout  nd_aib9_ch4_x0y0, 
	inout  nd_aib8_ch4_x0y0, 
	inout  nd_aib7_ch4_x0y0, 
	inout  nd_aib6_ch4_x0y0, 
	inout  nd_aib5_ch4_x0y0, 
	inout  nd_aib4_ch4_x0y0, 
	inout  nd_aib3_ch4_x0y0, 
	inout  nd_aib2_ch4_x0y0, 
	inout  nd_aib1_ch4_x0y0, 
	inout  nd_aib0_ch4_x0y0, 
// ## START OF  ch5 ( ##
        inout [95:0] m0_ch5_aib,
 	inout  nd_aib95_ch5_x0y0, 
	inout  nd_aib94_ch5_x0y0, 
	inout  nd_aib93_ch5_x0y0, 
	inout  nd_aib92_ch5_x0y0, 
	inout  nd_aib91_ch5_x0y0, 
	inout  nd_aib90_ch5_x0y0, 
	inout  nd_aib89_ch5_x0y0, 
	inout  nd_aib88_ch5_x0y0, 
	inout  nd_aib87_ch5_x0y0, 
	inout  nd_aib86_ch5_x0y0, 
	inout  nd_aib85_ch5_x0y0, 
	inout  nd_aib84_ch5_x0y0, 
	inout  nd_aib83_ch5_x0y0, 
	inout  nd_aib82_ch5_x0y0, 
	inout  nd_aib81_ch5_x0y0, 
	inout  nd_aib80_ch5_x0y0, 
	inout  nd_aib79_ch5_x0y0, 
	inout  nd_aib78_ch5_x0y0, 
	inout  nd_aib77_ch5_x0y0, 
	inout  nd_aib76_ch5_x0y0, 
	inout  nd_aib75_ch5_x0y0, 
	inout  nd_aib74_ch5_x0y0, 
	inout  nd_aib73_ch5_x0y0, 
	inout  nd_aib72_ch5_x0y0, 
	inout  nd_aib71_ch5_x0y0, 
	inout  nd_aib70_ch5_x0y0, 
	inout  nd_aib69_ch5_x0y0, 
	inout  nd_aib68_ch5_x0y0, 
	inout  nd_aib67_ch5_x0y0, 
	inout  nd_aib66_ch5_x0y0, 
	inout  nd_aib65_ch5_x0y0, 
	inout  nd_aib64_ch5_x0y0, 
	inout  nd_aib63_ch5_x0y0, 
	inout  nd_aib62_ch5_x0y0, 
	inout  nd_aib61_ch5_x0y0, 
	inout  nd_aib60_ch5_x0y0, 
	inout  nd_aib59_ch5_x0y0, 
	inout  nd_aib58_ch5_x0y0, 
	inout  nd_aib57_ch5_x0y0, 
	inout  nd_aib56_ch5_x0y0, 
	inout  nd_aib55_ch5_x0y0, 
	inout  nd_aib54_ch5_x0y0, 
	inout  nd_aib53_ch5_x0y0, 
	inout  nd_aib52_ch5_x0y0, 
	inout  nd_aib51_ch5_x0y0, 
	inout  nd_aib50_ch5_x0y0, 
	inout  nd_aib49_ch5_x0y0, 
	inout  nd_aib48_ch5_x0y0, 
	inout  nd_aib47_ch5_x0y0, 
	inout  nd_aib46_ch5_x0y0, 
	inout  nd_aib45_ch5_x0y0, 
	inout  nd_aib44_ch5_x0y0, 
	inout  nd_aib43_ch5_x0y0, 
	inout  nd_aib42_ch5_x0y0, 
	inout  nd_aib41_ch5_x0y0, 
	inout  nd_aib40_ch5_x0y0, 
	inout  nd_aib39_ch5_x0y0, 
	inout  nd_aib38_ch5_x0y0, 
	inout  nd_aib37_ch5_x0y0, 
	inout  nd_aib36_ch5_x0y0, 
	inout  nd_aib35_ch5_x0y0, 
	inout  nd_aib34_ch5_x0y0, 
	inout  nd_aib33_ch5_x0y0, 
	inout  nd_aib32_ch5_x0y0, 
	inout  nd_aib31_ch5_x0y0, 
	inout  nd_aib30_ch5_x0y0, 
	inout  nd_aib29_ch5_x0y0, 
	inout  nd_aib28_ch5_x0y0, 
	inout  nd_aib27_ch5_x0y0, 
	inout  nd_aib26_ch5_x0y0, 
	inout  nd_aib25_ch5_x0y0, 
	inout  nd_aib24_ch5_x0y0, 
	inout  nd_aib23_ch5_x0y0, 
	inout  nd_aib22_ch5_x0y0, 
	inout  nd_aib21_ch5_x0y0, 
	inout  nd_aib20_ch5_x0y0, 
	inout  nd_aib19_ch5_x0y0, 
	inout  nd_aib18_ch5_x0y0, 
	inout  nd_aib17_ch5_x0y0, 
	inout  nd_aib16_ch5_x0y0, 
	inout  nd_aib15_ch5_x0y0, 
	inout  nd_aib14_ch5_x0y0, 
	inout  nd_aib13_ch5_x0y0, 
	inout  nd_aib12_ch5_x0y0, 
	inout  nd_aib11_ch5_x0y0, 
	inout  nd_aib10_ch5_x0y0, 
	inout  nd_aib9_ch5_x0y0, 
	inout  nd_aib8_ch5_x0y0, 
	inout  nd_aib7_ch5_x0y0, 
	inout  nd_aib6_ch5_x0y0, 
	inout  nd_aib5_ch5_x0y0, 
	inout  nd_aib4_ch5_x0y0, 
	inout  nd_aib3_ch5_x0y0, 
	inout  nd_aib2_ch5_x0y0, 
	inout  nd_aib1_ch5_x0y0, 
	inout  nd_aib0_ch5_x0y0, 
// ## START OF  ch6 ( ##
        inout [95:0] m1_ch0_aib,
 	inout  nd_aib95_ch0_x0y1, 
	inout  nd_aib94_ch0_x0y1, 
	inout  nd_aib93_ch0_x0y1, 
	inout  nd_aib92_ch0_x0y1, 
	inout  nd_aib91_ch0_x0y1, 
	inout  nd_aib90_ch0_x0y1, 
	inout  nd_aib89_ch0_x0y1, 
	inout  nd_aib88_ch0_x0y1, 
	inout  nd_aib87_ch0_x0y1, 
	inout  nd_aib86_ch0_x0y1, 
	inout  nd_aib85_ch0_x0y1, 
	inout  nd_aib84_ch0_x0y1, 
	inout  nd_aib83_ch0_x0y1, 
	inout  nd_aib82_ch0_x0y1, 
	inout  nd_aib81_ch0_x0y1, 
	inout  nd_aib80_ch0_x0y1, 
	inout  nd_aib79_ch0_x0y1, 
	inout  nd_aib78_ch0_x0y1, 
	inout  nd_aib77_ch0_x0y1, 
	inout  nd_aib76_ch0_x0y1, 
	inout  nd_aib75_ch0_x0y1, 
	inout  nd_aib74_ch0_x0y1, 
	inout  nd_aib73_ch0_x0y1, 
	inout  nd_aib72_ch0_x0y1, 
	inout  nd_aib71_ch0_x0y1, 
	inout  nd_aib70_ch0_x0y1, 
	inout  nd_aib69_ch0_x0y1, 
	inout  nd_aib68_ch0_x0y1, 
	inout  nd_aib67_ch0_x0y1, 
	inout  nd_aib66_ch0_x0y1, 
	inout  nd_aib65_ch0_x0y1, 
	inout  nd_aib64_ch0_x0y1, 
	inout  nd_aib63_ch0_x0y1, 
	inout  nd_aib62_ch0_x0y1, 
	inout  nd_aib61_ch0_x0y1, 
	inout  nd_aib60_ch0_x0y1, 
	inout  nd_aib59_ch0_x0y1, 
	inout  nd_aib58_ch0_x0y1, 
	inout  nd_aib57_ch0_x0y1, 
	inout  nd_aib56_ch0_x0y1, 
	inout  nd_aib55_ch0_x0y1, 
	inout  nd_aib54_ch0_x0y1, 
	inout  nd_aib53_ch0_x0y1, 
	inout  nd_aib52_ch0_x0y1, 
	inout  nd_aib51_ch0_x0y1, 
	inout  nd_aib50_ch0_x0y1, 
	inout  nd_aib49_ch0_x0y1, 
	inout  nd_aib48_ch0_x0y1, 
	inout  nd_aib47_ch0_x0y1, 
	inout  nd_aib46_ch0_x0y1, 
	inout  nd_aib45_ch0_x0y1, 
	inout  nd_aib44_ch0_x0y1, 
	inout  nd_aib43_ch0_x0y1, 
	inout  nd_aib42_ch0_x0y1, 
	inout  nd_aib41_ch0_x0y1, 
	inout  nd_aib40_ch0_x0y1, 
	inout  nd_aib39_ch0_x0y1, 
	inout  nd_aib38_ch0_x0y1, 
	inout  nd_aib37_ch0_x0y1, 
	inout  nd_aib36_ch0_x0y1, 
	inout  nd_aib35_ch0_x0y1, 
	inout  nd_aib34_ch0_x0y1, 
	inout  nd_aib33_ch0_x0y1, 
	inout  nd_aib32_ch0_x0y1, 
	inout  nd_aib31_ch0_x0y1, 
	inout  nd_aib30_ch0_x0y1, 
	inout  nd_aib29_ch0_x0y1, 
	inout  nd_aib28_ch0_x0y1, 
	inout  nd_aib27_ch0_x0y1, 
	inout  nd_aib26_ch0_x0y1, 
	inout  nd_aib25_ch0_x0y1, 
	inout  nd_aib24_ch0_x0y1, 
	inout  nd_aib23_ch0_x0y1, 
	inout  nd_aib22_ch0_x0y1, 
	inout  nd_aib21_ch0_x0y1, 
	inout  nd_aib20_ch0_x0y1, 
	inout  nd_aib19_ch0_x0y1, 
	inout  nd_aib18_ch0_x0y1, 
	inout  nd_aib17_ch0_x0y1, 
	inout  nd_aib16_ch0_x0y1, 
	inout  nd_aib15_ch0_x0y1, 
	inout  nd_aib14_ch0_x0y1, 
	inout  nd_aib13_ch0_x0y1, 
	inout  nd_aib12_ch0_x0y1, 
	inout  nd_aib11_ch0_x0y1, 
	inout  nd_aib10_ch0_x0y1, 
	inout  nd_aib9_ch0_x0y1, 
	inout  nd_aib8_ch0_x0y1, 
	inout  nd_aib7_ch0_x0y1, 
	inout  nd_aib6_ch0_x0y1, 
	inout  nd_aib5_ch0_x0y1, 
	inout  nd_aib4_ch0_x0y1, 
	inout  nd_aib3_ch0_x0y1, 
	inout  nd_aib2_ch0_x0y1, 
	inout  nd_aib1_ch0_x0y1, 
	inout  nd_aib0_ch0_x0y1, 
// ## START OF  ch7 ( ##
        inout [95:0] m1_ch1_aib,
 	inout  nd_aib95_ch1_x0y1, 
	inout  nd_aib94_ch1_x0y1, 
	inout  nd_aib93_ch1_x0y1, 
	inout  nd_aib92_ch1_x0y1, 
	inout  nd_aib91_ch1_x0y1, 
	inout  nd_aib90_ch1_x0y1, 
	inout  nd_aib89_ch1_x0y1, 
	inout  nd_aib88_ch1_x0y1, 
	inout  nd_aib87_ch1_x0y1, 
	inout  nd_aib86_ch1_x0y1, 
	inout  nd_aib85_ch1_x0y1, 
	inout  nd_aib84_ch1_x0y1, 
	inout  nd_aib83_ch1_x0y1, 
	inout  nd_aib82_ch1_x0y1, 
	inout  nd_aib81_ch1_x0y1, 
	inout  nd_aib80_ch1_x0y1, 
	inout  nd_aib79_ch1_x0y1, 
	inout  nd_aib78_ch1_x0y1, 
	inout  nd_aib77_ch1_x0y1, 
	inout  nd_aib76_ch1_x0y1, 
	inout  nd_aib75_ch1_x0y1, 
	inout  nd_aib74_ch1_x0y1, 
	inout  nd_aib73_ch1_x0y1, 
	inout  nd_aib72_ch1_x0y1, 
	inout  nd_aib71_ch1_x0y1, 
	inout  nd_aib70_ch1_x0y1, 
	inout  nd_aib69_ch1_x0y1, 
	inout  nd_aib68_ch1_x0y1, 
	inout  nd_aib67_ch1_x0y1, 
	inout  nd_aib66_ch1_x0y1, 
	inout  nd_aib65_ch1_x0y1, 
	inout  nd_aib64_ch1_x0y1, 
	inout  nd_aib63_ch1_x0y1, 
	inout  nd_aib62_ch1_x0y1, 
	inout  nd_aib61_ch1_x0y1, 
	inout  nd_aib60_ch1_x0y1, 
	inout  nd_aib59_ch1_x0y1, 
	inout  nd_aib58_ch1_x0y1, 
	inout  nd_aib57_ch1_x0y1, 
	inout  nd_aib56_ch1_x0y1, 
	inout  nd_aib55_ch1_x0y1, 
	inout  nd_aib54_ch1_x0y1, 
	inout  nd_aib53_ch1_x0y1, 
	inout  nd_aib52_ch1_x0y1, 
	inout  nd_aib51_ch1_x0y1, 
	inout  nd_aib50_ch1_x0y1, 
	inout  nd_aib49_ch1_x0y1, 
	inout  nd_aib48_ch1_x0y1, 
	inout  nd_aib47_ch1_x0y1, 
	inout  nd_aib46_ch1_x0y1, 
	inout  nd_aib45_ch1_x0y1, 
	inout  nd_aib44_ch1_x0y1, 
	inout  nd_aib43_ch1_x0y1, 
	inout  nd_aib42_ch1_x0y1, 
	inout  nd_aib41_ch1_x0y1, 
	inout  nd_aib40_ch1_x0y1, 
	inout  nd_aib39_ch1_x0y1, 
	inout  nd_aib38_ch1_x0y1, 
	inout  nd_aib37_ch1_x0y1, 
	inout  nd_aib36_ch1_x0y1, 
	inout  nd_aib35_ch1_x0y1, 
	inout  nd_aib34_ch1_x0y1, 
	inout  nd_aib33_ch1_x0y1, 
	inout  nd_aib32_ch1_x0y1, 
	inout  nd_aib31_ch1_x0y1, 
	inout  nd_aib30_ch1_x0y1, 
	inout  nd_aib29_ch1_x0y1, 
	inout  nd_aib28_ch1_x0y1, 
	inout  nd_aib27_ch1_x0y1, 
	inout  nd_aib26_ch1_x0y1, 
	inout  nd_aib25_ch1_x0y1, 
	inout  nd_aib24_ch1_x0y1, 
	inout  nd_aib23_ch1_x0y1, 
	inout  nd_aib22_ch1_x0y1, 
	inout  nd_aib21_ch1_x0y1, 
	inout  nd_aib20_ch1_x0y1, 
	inout  nd_aib19_ch1_x0y1, 
	inout  nd_aib18_ch1_x0y1, 
	inout  nd_aib17_ch1_x0y1, 
	inout  nd_aib16_ch1_x0y1, 
	inout  nd_aib15_ch1_x0y1, 
	inout  nd_aib14_ch1_x0y1, 
	inout  nd_aib13_ch1_x0y1, 
	inout  nd_aib12_ch1_x0y1, 
	inout  nd_aib11_ch1_x0y1, 
	inout  nd_aib10_ch1_x0y1, 
	inout  nd_aib9_ch1_x0y1, 
	inout  nd_aib8_ch1_x0y1, 
	inout  nd_aib7_ch1_x0y1, 
	inout  nd_aib6_ch1_x0y1, 
	inout  nd_aib5_ch1_x0y1, 
	inout  nd_aib4_ch1_x0y1, 
	inout  nd_aib3_ch1_x0y1, 
	inout  nd_aib2_ch1_x0y1, 
	inout  nd_aib1_ch1_x0y1, 
	inout  nd_aib0_ch1_x0y1, 
// ## START OF  ch8 ( ##
        inout [95:0] m1_ch2_aib,
 	inout  nd_aib95_ch2_x0y1, 
	inout  nd_aib94_ch2_x0y1, 
	inout  nd_aib93_ch2_x0y1, 
	inout  nd_aib92_ch2_x0y1, 
	inout  nd_aib91_ch2_x0y1, 
	inout  nd_aib90_ch2_x0y1, 
	inout  nd_aib89_ch2_x0y1, 
	inout  nd_aib88_ch2_x0y1, 
	inout  nd_aib87_ch2_x0y1, 
	inout  nd_aib86_ch2_x0y1, 
	inout  nd_aib85_ch2_x0y1, 
	inout  nd_aib84_ch2_x0y1, 
	inout  nd_aib83_ch2_x0y1, 
	inout  nd_aib82_ch2_x0y1, 
	inout  nd_aib81_ch2_x0y1, 
	inout  nd_aib80_ch2_x0y1, 
	inout  nd_aib79_ch2_x0y1, 
	inout  nd_aib78_ch2_x0y1, 
	inout  nd_aib77_ch2_x0y1, 
	inout  nd_aib76_ch2_x0y1, 
	inout  nd_aib75_ch2_x0y1, 
	inout  nd_aib74_ch2_x0y1, 
	inout  nd_aib73_ch2_x0y1, 
	inout  nd_aib72_ch2_x0y1, 
	inout  nd_aib71_ch2_x0y1, 
	inout  nd_aib70_ch2_x0y1, 
	inout  nd_aib69_ch2_x0y1, 
	inout  nd_aib68_ch2_x0y1, 
	inout  nd_aib67_ch2_x0y1, 
	inout  nd_aib66_ch2_x0y1, 
	inout  nd_aib65_ch2_x0y1, 
	inout  nd_aib64_ch2_x0y1, 
	inout  nd_aib63_ch2_x0y1, 
	inout  nd_aib62_ch2_x0y1, 
	inout  nd_aib61_ch2_x0y1, 
	inout  nd_aib60_ch2_x0y1, 
	inout  nd_aib59_ch2_x0y1, 
	inout  nd_aib58_ch2_x0y1, 
	inout  nd_aib57_ch2_x0y1, 
	inout  nd_aib56_ch2_x0y1, 
	inout  nd_aib55_ch2_x0y1, 
	inout  nd_aib54_ch2_x0y1, 
	inout  nd_aib53_ch2_x0y1, 
	inout  nd_aib52_ch2_x0y1, 
	inout  nd_aib51_ch2_x0y1, 
	inout  nd_aib50_ch2_x0y1, 
	inout  nd_aib49_ch2_x0y1, 
	inout  nd_aib48_ch2_x0y1, 
	inout  nd_aib47_ch2_x0y1, 
	inout  nd_aib46_ch2_x0y1, 
	inout  nd_aib45_ch2_x0y1, 
	inout  nd_aib44_ch2_x0y1, 
	inout  nd_aib43_ch2_x0y1, 
	inout  nd_aib42_ch2_x0y1, 
	inout  nd_aib41_ch2_x0y1, 
	inout  nd_aib40_ch2_x0y1, 
	inout  nd_aib39_ch2_x0y1, 
	inout  nd_aib38_ch2_x0y1, 
	inout  nd_aib37_ch2_x0y1, 
	inout  nd_aib36_ch2_x0y1, 
	inout  nd_aib35_ch2_x0y1, 
	inout  nd_aib34_ch2_x0y1, 
	inout  nd_aib33_ch2_x0y1, 
	inout  nd_aib32_ch2_x0y1, 
	inout  nd_aib31_ch2_x0y1, 
	inout  nd_aib30_ch2_x0y1, 
	inout  nd_aib29_ch2_x0y1, 
	inout  nd_aib28_ch2_x0y1, 
	inout  nd_aib27_ch2_x0y1, 
	inout  nd_aib26_ch2_x0y1, 
	inout  nd_aib25_ch2_x0y1, 
	inout  nd_aib24_ch2_x0y1, 
	inout  nd_aib23_ch2_x0y1, 
	inout  nd_aib22_ch2_x0y1, 
	inout  nd_aib21_ch2_x0y1, 
	inout  nd_aib20_ch2_x0y1, 
	inout  nd_aib19_ch2_x0y1, 
	inout  nd_aib18_ch2_x0y1, 
	inout  nd_aib17_ch2_x0y1, 
	inout  nd_aib16_ch2_x0y1, 
	inout  nd_aib15_ch2_x0y1, 
	inout  nd_aib14_ch2_x0y1, 
	inout  nd_aib13_ch2_x0y1, 
	inout  nd_aib12_ch2_x0y1, 
	inout  nd_aib11_ch2_x0y1, 
	inout  nd_aib10_ch2_x0y1, 
	inout  nd_aib9_ch2_x0y1, 
	inout  nd_aib8_ch2_x0y1, 
	inout  nd_aib7_ch2_x0y1, 
	inout  nd_aib6_ch2_x0y1, 
	inout  nd_aib5_ch2_x0y1, 
	inout  nd_aib4_ch2_x0y1, 
	inout  nd_aib3_ch2_x0y1, 
	inout  nd_aib2_ch2_x0y1, 
	inout  nd_aib1_ch2_x0y1, 
	inout  nd_aib0_ch2_x0y1, 
// ## START OF  ch9 ( ##
        inout [95:0] m1_ch3_aib,
 	inout  nd_aib95_ch3_x0y1, 
	inout  nd_aib94_ch3_x0y1, 
	inout  nd_aib93_ch3_x0y1, 
	inout  nd_aib92_ch3_x0y1, 
	inout  nd_aib91_ch3_x0y1, 
	inout  nd_aib90_ch3_x0y1, 
	inout  nd_aib89_ch3_x0y1, 
	inout  nd_aib88_ch3_x0y1, 
	inout  nd_aib87_ch3_x0y1, 
	inout  nd_aib86_ch3_x0y1, 
	inout  nd_aib85_ch3_x0y1, 
	inout  nd_aib84_ch3_x0y1, 
	inout  nd_aib83_ch3_x0y1, 
	inout  nd_aib82_ch3_x0y1, 
	inout  nd_aib81_ch3_x0y1, 
	inout  nd_aib80_ch3_x0y1, 
	inout  nd_aib79_ch3_x0y1, 
	inout  nd_aib78_ch3_x0y1, 
	inout  nd_aib77_ch3_x0y1, 
	inout  nd_aib76_ch3_x0y1, 
	inout  nd_aib75_ch3_x0y1, 
	inout  nd_aib74_ch3_x0y1, 
	inout  nd_aib73_ch3_x0y1, 
	inout  nd_aib72_ch3_x0y1, 
	inout  nd_aib71_ch3_x0y1, 
	inout  nd_aib70_ch3_x0y1, 
	inout  nd_aib69_ch3_x0y1, 
	inout  nd_aib68_ch3_x0y1, 
	inout  nd_aib67_ch3_x0y1, 
	inout  nd_aib66_ch3_x0y1, 
	inout  nd_aib65_ch3_x0y1, 
	inout  nd_aib64_ch3_x0y1, 
	inout  nd_aib63_ch3_x0y1, 
	inout  nd_aib62_ch3_x0y1, 
	inout  nd_aib61_ch3_x0y1, 
	inout  nd_aib60_ch3_x0y1, 
	inout  nd_aib59_ch3_x0y1, 
	inout  nd_aib58_ch3_x0y1, 
	inout  nd_aib57_ch3_x0y1, 
	inout  nd_aib56_ch3_x0y1, 
	inout  nd_aib55_ch3_x0y1, 
	inout  nd_aib54_ch3_x0y1, 
	inout  nd_aib53_ch3_x0y1, 
	inout  nd_aib52_ch3_x0y1, 
	inout  nd_aib51_ch3_x0y1, 
	inout  nd_aib50_ch3_x0y1, 
	inout  nd_aib49_ch3_x0y1, 
	inout  nd_aib48_ch3_x0y1, 
	inout  nd_aib47_ch3_x0y1, 
	inout  nd_aib46_ch3_x0y1, 
	inout  nd_aib45_ch3_x0y1, 
	inout  nd_aib44_ch3_x0y1, 
	inout  nd_aib43_ch3_x0y1, 
	inout  nd_aib42_ch3_x0y1, 
	inout  nd_aib41_ch3_x0y1, 
	inout  nd_aib40_ch3_x0y1, 
	inout  nd_aib39_ch3_x0y1, 
	inout  nd_aib38_ch3_x0y1, 
	inout  nd_aib37_ch3_x0y1, 
	inout  nd_aib36_ch3_x0y1, 
	inout  nd_aib35_ch3_x0y1, 
	inout  nd_aib34_ch3_x0y1, 
	inout  nd_aib33_ch3_x0y1, 
	inout  nd_aib32_ch3_x0y1, 
	inout  nd_aib31_ch3_x0y1, 
	inout  nd_aib30_ch3_x0y1, 
	inout  nd_aib29_ch3_x0y1, 
	inout  nd_aib28_ch3_x0y1, 
	inout  nd_aib27_ch3_x0y1, 
	inout  nd_aib26_ch3_x0y1, 
	inout  nd_aib25_ch3_x0y1, 
	inout  nd_aib24_ch3_x0y1, 
	inout  nd_aib23_ch3_x0y1, 
	inout  nd_aib22_ch3_x0y1, 
	inout  nd_aib21_ch3_x0y1, 
	inout  nd_aib20_ch3_x0y1, 
	inout  nd_aib19_ch3_x0y1, 
	inout  nd_aib18_ch3_x0y1, 
	inout  nd_aib17_ch3_x0y1, 
	inout  nd_aib16_ch3_x0y1, 
	inout  nd_aib15_ch3_x0y1, 
	inout  nd_aib14_ch3_x0y1, 
	inout  nd_aib13_ch3_x0y1, 
	inout  nd_aib12_ch3_x0y1, 
	inout  nd_aib11_ch3_x0y1, 
	inout  nd_aib10_ch3_x0y1, 
	inout  nd_aib9_ch3_x0y1, 
	inout  nd_aib8_ch3_x0y1, 
	inout  nd_aib7_ch3_x0y1, 
	inout  nd_aib6_ch3_x0y1, 
	inout  nd_aib5_ch3_x0y1, 
	inout  nd_aib4_ch3_x0y1, 
	inout  nd_aib3_ch3_x0y1, 
	inout  nd_aib2_ch3_x0y1, 
	inout  nd_aib1_ch3_x0y1, 
	inout  nd_aib0_ch3_x0y1, 
// ## START OF  ch10 ( ##
        inout [95:0] m1_ch4_aib,
 	inout  nd_aib95_ch4_x0y1, 
	inout  nd_aib94_ch4_x0y1, 
	inout  nd_aib93_ch4_x0y1, 
	inout  nd_aib92_ch4_x0y1, 
	inout  nd_aib91_ch4_x0y1, 
	inout  nd_aib90_ch4_x0y1, 
	inout  nd_aib89_ch4_x0y1, 
	inout  nd_aib88_ch4_x0y1, 
	inout  nd_aib87_ch4_x0y1, 
	inout  nd_aib86_ch4_x0y1, 
	inout  nd_aib85_ch4_x0y1, 
	inout  nd_aib84_ch4_x0y1, 
	inout  nd_aib83_ch4_x0y1, 
	inout  nd_aib82_ch4_x0y1, 
	inout  nd_aib81_ch4_x0y1, 
	inout  nd_aib80_ch4_x0y1, 
	inout  nd_aib79_ch4_x0y1, 
	inout  nd_aib78_ch4_x0y1, 
	inout  nd_aib77_ch4_x0y1, 
	inout  nd_aib76_ch4_x0y1, 
	inout  nd_aib75_ch4_x0y1, 
	inout  nd_aib74_ch4_x0y1, 
	inout  nd_aib73_ch4_x0y1, 
	inout  nd_aib72_ch4_x0y1, 
	inout  nd_aib71_ch4_x0y1, 
	inout  nd_aib70_ch4_x0y1, 
	inout  nd_aib69_ch4_x0y1, 
	inout  nd_aib68_ch4_x0y1, 
	inout  nd_aib67_ch4_x0y1, 
	inout  nd_aib66_ch4_x0y1, 
	inout  nd_aib65_ch4_x0y1, 
	inout  nd_aib64_ch4_x0y1, 
	inout  nd_aib63_ch4_x0y1, 
	inout  nd_aib62_ch4_x0y1, 
	inout  nd_aib61_ch4_x0y1, 
	inout  nd_aib60_ch4_x0y1, 
	inout  nd_aib59_ch4_x0y1, 
	inout  nd_aib58_ch4_x0y1, 
	inout  nd_aib57_ch4_x0y1, 
	inout  nd_aib56_ch4_x0y1, 
	inout  nd_aib55_ch4_x0y1, 
	inout  nd_aib54_ch4_x0y1, 
	inout  nd_aib53_ch4_x0y1, 
	inout  nd_aib52_ch4_x0y1, 
	inout  nd_aib51_ch4_x0y1, 
	inout  nd_aib50_ch4_x0y1, 
	inout  nd_aib49_ch4_x0y1, 
	inout  nd_aib48_ch4_x0y1, 
	inout  nd_aib47_ch4_x0y1, 
	inout  nd_aib46_ch4_x0y1, 
	inout  nd_aib45_ch4_x0y1, 
	inout  nd_aib44_ch4_x0y1, 
	inout  nd_aib43_ch4_x0y1, 
	inout  nd_aib42_ch4_x0y1, 
	inout  nd_aib41_ch4_x0y1, 
	inout  nd_aib40_ch4_x0y1, 
	inout  nd_aib39_ch4_x0y1, 
	inout  nd_aib38_ch4_x0y1, 
	inout  nd_aib37_ch4_x0y1, 
	inout  nd_aib36_ch4_x0y1, 
	inout  nd_aib35_ch4_x0y1, 
	inout  nd_aib34_ch4_x0y1, 
	inout  nd_aib33_ch4_x0y1, 
	inout  nd_aib32_ch4_x0y1, 
	inout  nd_aib31_ch4_x0y1, 
	inout  nd_aib30_ch4_x0y1, 
	inout  nd_aib29_ch4_x0y1, 
	inout  nd_aib28_ch4_x0y1, 
	inout  nd_aib27_ch4_x0y1, 
	inout  nd_aib26_ch4_x0y1, 
	inout  nd_aib25_ch4_x0y1, 
	inout  nd_aib24_ch4_x0y1, 
	inout  nd_aib23_ch4_x0y1, 
	inout  nd_aib22_ch4_x0y1, 
	inout  nd_aib21_ch4_x0y1, 
	inout  nd_aib20_ch4_x0y1, 
	inout  nd_aib19_ch4_x0y1, 
	inout  nd_aib18_ch4_x0y1, 
	inout  nd_aib17_ch4_x0y1, 
	inout  nd_aib16_ch4_x0y1, 
	inout  nd_aib15_ch4_x0y1, 
	inout  nd_aib14_ch4_x0y1, 
	inout  nd_aib13_ch4_x0y1, 
	inout  nd_aib12_ch4_x0y1, 
	inout  nd_aib11_ch4_x0y1, 
	inout  nd_aib10_ch4_x0y1, 
	inout  nd_aib9_ch4_x0y1, 
	inout  nd_aib8_ch4_x0y1, 
	inout  nd_aib7_ch4_x0y1, 
	inout  nd_aib6_ch4_x0y1, 
	inout  nd_aib5_ch4_x0y1, 
	inout  nd_aib4_ch4_x0y1, 
	inout  nd_aib3_ch4_x0y1, 
	inout  nd_aib2_ch4_x0y1, 
	inout  nd_aib1_ch4_x0y1, 
	inout  nd_aib0_ch4_x0y1, 
// ## START OF  ch11 ( ##
        inout [95:0] m1_ch5_aib,
 	inout  nd_aib95_ch5_x0y1, 
	inout  nd_aib94_ch5_x0y1, 
	inout  nd_aib93_ch5_x0y1, 
	inout  nd_aib92_ch5_x0y1, 
	inout  nd_aib91_ch5_x0y1, 
	inout  nd_aib90_ch5_x0y1, 
	inout  nd_aib89_ch5_x0y1, 
	inout  nd_aib88_ch5_x0y1, 
	inout  nd_aib87_ch5_x0y1, 
	inout  nd_aib86_ch5_x0y1, 
	inout  nd_aib85_ch5_x0y1, 
	inout  nd_aib84_ch5_x0y1, 
	inout  nd_aib83_ch5_x0y1, 
	inout  nd_aib82_ch5_x0y1, 
	inout  nd_aib81_ch5_x0y1, 
	inout  nd_aib80_ch5_x0y1, 
	inout  nd_aib79_ch5_x0y1, 
	inout  nd_aib78_ch5_x0y1, 
	inout  nd_aib77_ch5_x0y1, 
	inout  nd_aib76_ch5_x0y1, 
	inout  nd_aib75_ch5_x0y1, 
	inout  nd_aib74_ch5_x0y1, 
	inout  nd_aib73_ch5_x0y1, 
	inout  nd_aib72_ch5_x0y1, 
	inout  nd_aib71_ch5_x0y1, 
	inout  nd_aib70_ch5_x0y1, 
	inout  nd_aib69_ch5_x0y1, 
	inout  nd_aib68_ch5_x0y1, 
	inout  nd_aib67_ch5_x0y1, 
	inout  nd_aib66_ch5_x0y1, 
	inout  nd_aib65_ch5_x0y1, 
	inout  nd_aib64_ch5_x0y1, 
	inout  nd_aib63_ch5_x0y1, 
	inout  nd_aib62_ch5_x0y1, 
	inout  nd_aib61_ch5_x0y1, 
	inout  nd_aib60_ch5_x0y1, 
	inout  nd_aib59_ch5_x0y1, 
	inout  nd_aib58_ch5_x0y1, 
	inout  nd_aib57_ch5_x0y1, 
	inout  nd_aib56_ch5_x0y1, 
	inout  nd_aib55_ch5_x0y1, 
	inout  nd_aib54_ch5_x0y1, 
	inout  nd_aib53_ch5_x0y1, 
	inout  nd_aib52_ch5_x0y1, 
	inout  nd_aib51_ch5_x0y1, 
	inout  nd_aib50_ch5_x0y1, 
	inout  nd_aib49_ch5_x0y1, 
	inout  nd_aib48_ch5_x0y1, 
	inout  nd_aib47_ch5_x0y1, 
	inout  nd_aib46_ch5_x0y1, 
	inout  nd_aib45_ch5_x0y1, 
	inout  nd_aib44_ch5_x0y1, 
	inout  nd_aib43_ch5_x0y1, 
	inout  nd_aib42_ch5_x0y1, 
	inout  nd_aib41_ch5_x0y1, 
	inout  nd_aib40_ch5_x0y1, 
	inout  nd_aib39_ch5_x0y1, 
	inout  nd_aib38_ch5_x0y1, 
	inout  nd_aib37_ch5_x0y1, 
	inout  nd_aib36_ch5_x0y1, 
	inout  nd_aib35_ch5_x0y1, 
	inout  nd_aib34_ch5_x0y1, 
	inout  nd_aib33_ch5_x0y1, 
	inout  nd_aib32_ch5_x0y1, 
	inout  nd_aib31_ch5_x0y1, 
	inout  nd_aib30_ch5_x0y1, 
	inout  nd_aib29_ch5_x0y1, 
	inout  nd_aib28_ch5_x0y1, 
	inout  nd_aib27_ch5_x0y1, 
	inout  nd_aib26_ch5_x0y1, 
	inout  nd_aib25_ch5_x0y1, 
	inout  nd_aib24_ch5_x0y1, 
	inout  nd_aib23_ch5_x0y1, 
	inout  nd_aib22_ch5_x0y1, 
	inout  nd_aib21_ch5_x0y1, 
	inout  nd_aib20_ch5_x0y1, 
	inout  nd_aib19_ch5_x0y1, 
	inout  nd_aib18_ch5_x0y1, 
	inout  nd_aib17_ch5_x0y1, 
	inout  nd_aib16_ch5_x0y1, 
	inout  nd_aib15_ch5_x0y1, 
	inout  nd_aib14_ch5_x0y1, 
	inout  nd_aib13_ch5_x0y1, 
	inout  nd_aib12_ch5_x0y1, 
	inout  nd_aib11_ch5_x0y1, 
	inout  nd_aib10_ch5_x0y1, 
	inout  nd_aib9_ch5_x0y1, 
	inout  nd_aib8_ch5_x0y1, 
	inout  nd_aib7_ch5_x0y1, 
	inout  nd_aib6_ch5_x0y1, 
	inout  nd_aib5_ch5_x0y1, 
	inout  nd_aib4_ch5_x0y1, 
	inout  nd_aib3_ch5_x0y1, 
	inout  nd_aib2_ch5_x0y1, 
	inout  nd_aib1_ch5_x0y1, 
	inout  nd_aib0_ch5_x0y1, 
// ## START OF ch12 ( ##
        inout [95:0] m2_ch0_aib,
 	inout  nd_aib95_ch0_x0y2, 
	inout  nd_aib94_ch0_x0y2, 
	inout  nd_aib93_ch0_x0y2, 
	inout  nd_aib92_ch0_x0y2, 
	inout  nd_aib91_ch0_x0y2, 
	inout  nd_aib90_ch0_x0y2, 
	inout  nd_aib89_ch0_x0y2, 
	inout  nd_aib88_ch0_x0y2, 
	inout  nd_aib87_ch0_x0y2, 
	inout  nd_aib86_ch0_x0y2, 
	inout  nd_aib85_ch0_x0y2, 
	inout  nd_aib84_ch0_x0y2, 
	inout  nd_aib83_ch0_x0y2, 
	inout  nd_aib82_ch0_x0y2, 
	inout  nd_aib81_ch0_x0y2, 
	inout  nd_aib80_ch0_x0y2, 
	inout  nd_aib79_ch0_x0y2, 
	inout  nd_aib78_ch0_x0y2, 
	inout  nd_aib77_ch0_x0y2, 
	inout  nd_aib76_ch0_x0y2, 
	inout  nd_aib75_ch0_x0y2, 
	inout  nd_aib74_ch0_x0y2, 
	inout  nd_aib73_ch0_x0y2, 
	inout  nd_aib72_ch0_x0y2, 
	inout  nd_aib71_ch0_x0y2, 
	inout  nd_aib70_ch0_x0y2, 
	inout  nd_aib69_ch0_x0y2, 
	inout  nd_aib68_ch0_x0y2, 
	inout  nd_aib67_ch0_x0y2, 
	inout  nd_aib66_ch0_x0y2, 
	inout  nd_aib65_ch0_x0y2, 
	inout  nd_aib64_ch0_x0y2, 
	inout  nd_aib63_ch0_x0y2, 
	inout  nd_aib62_ch0_x0y2, 
	inout  nd_aib61_ch0_x0y2, 
	inout  nd_aib60_ch0_x0y2, 
	inout  nd_aib59_ch0_x0y2, 
	inout  nd_aib58_ch0_x0y2, 
	inout  nd_aib57_ch0_x0y2, 
	inout  nd_aib56_ch0_x0y2, 
	inout  nd_aib55_ch0_x0y2, 
	inout  nd_aib54_ch0_x0y2, 
	inout  nd_aib53_ch0_x0y2, 
	inout  nd_aib52_ch0_x0y2, 
	inout  nd_aib51_ch0_x0y2, 
	inout  nd_aib50_ch0_x0y2, 
	inout  nd_aib49_ch0_x0y2, 
	inout  nd_aib48_ch0_x0y2, 
	inout  nd_aib47_ch0_x0y2, 
	inout  nd_aib46_ch0_x0y2, 
	inout  nd_aib45_ch0_x0y2, 
	inout  nd_aib44_ch0_x0y2, 
	inout  nd_aib43_ch0_x0y2, 
	inout  nd_aib42_ch0_x0y2, 
	inout  nd_aib41_ch0_x0y2, 
	inout  nd_aib40_ch0_x0y2, 
	inout  nd_aib39_ch0_x0y2, 
	inout  nd_aib38_ch0_x0y2, 
	inout  nd_aib37_ch0_x0y2, 
	inout  nd_aib36_ch0_x0y2, 
	inout  nd_aib35_ch0_x0y2, 
	inout  nd_aib34_ch0_x0y2, 
	inout  nd_aib33_ch0_x0y2, 
	inout  nd_aib32_ch0_x0y2, 
	inout  nd_aib31_ch0_x0y2, 
	inout  nd_aib30_ch0_x0y2, 
	inout  nd_aib29_ch0_x0y2, 
	inout  nd_aib28_ch0_x0y2, 
	inout  nd_aib27_ch0_x0y2, 
	inout  nd_aib26_ch0_x0y2, 
	inout  nd_aib25_ch0_x0y2, 
	inout  nd_aib24_ch0_x0y2, 
	inout  nd_aib23_ch0_x0y2, 
	inout  nd_aib22_ch0_x0y2, 
	inout  nd_aib21_ch0_x0y2, 
	inout  nd_aib20_ch0_x0y2, 
	inout  nd_aib19_ch0_x0y2, 
	inout  nd_aib18_ch0_x0y2, 
	inout  nd_aib17_ch0_x0y2, 
	inout  nd_aib16_ch0_x0y2, 
	inout  nd_aib15_ch0_x0y2, 
	inout  nd_aib14_ch0_x0y2, 
	inout  nd_aib13_ch0_x0y2, 
	inout  nd_aib12_ch0_x0y2, 
	inout  nd_aib11_ch0_x0y2, 
	inout  nd_aib10_ch0_x0y2, 
	inout  nd_aib9_ch0_x0y2, 
	inout  nd_aib8_ch0_x0y2, 
	inout  nd_aib7_ch0_x0y2, 
	inout  nd_aib6_ch0_x0y2, 
	inout  nd_aib5_ch0_x0y2, 
	inout  nd_aib4_ch0_x0y2, 
	inout  nd_aib3_ch0_x0y2, 
	inout  nd_aib2_ch0_x0y2, 
	inout  nd_aib1_ch0_x0y2, 
	inout  nd_aib0_ch0_x0y2, 
// ## START OF ch13 ( ##
        inout [95:0] m2_ch1_aib,
 	inout  nd_aib95_ch1_x0y2, 
	inout  nd_aib94_ch1_x0y2, 
	inout  nd_aib93_ch1_x0y2, 
	inout  nd_aib92_ch1_x0y2, 
	inout  nd_aib91_ch1_x0y2, 
	inout  nd_aib90_ch1_x0y2, 
	inout  nd_aib89_ch1_x0y2, 
	inout  nd_aib88_ch1_x0y2, 
	inout  nd_aib87_ch1_x0y2, 
	inout  nd_aib86_ch1_x0y2, 
	inout  nd_aib85_ch1_x0y2, 
	inout  nd_aib84_ch1_x0y2, 
	inout  nd_aib83_ch1_x0y2, 
	inout  nd_aib82_ch1_x0y2, 
	inout  nd_aib81_ch1_x0y2, 
	inout  nd_aib80_ch1_x0y2, 
	inout  nd_aib79_ch1_x0y2, 
	inout  nd_aib78_ch1_x0y2, 
	inout  nd_aib77_ch1_x0y2, 
	inout  nd_aib76_ch1_x0y2, 
	inout  nd_aib75_ch1_x0y2, 
	inout  nd_aib74_ch1_x0y2, 
	inout  nd_aib73_ch1_x0y2, 
	inout  nd_aib72_ch1_x0y2, 
	inout  nd_aib71_ch1_x0y2, 
	inout  nd_aib70_ch1_x0y2, 
	inout  nd_aib69_ch1_x0y2, 
	inout  nd_aib68_ch1_x0y2, 
	inout  nd_aib67_ch1_x0y2, 
	inout  nd_aib66_ch1_x0y2, 
	inout  nd_aib65_ch1_x0y2, 
	inout  nd_aib64_ch1_x0y2, 
	inout  nd_aib63_ch1_x0y2, 
	inout  nd_aib62_ch1_x0y2, 
	inout  nd_aib61_ch1_x0y2, 
	inout  nd_aib60_ch1_x0y2, 
	inout  nd_aib59_ch1_x0y2, 
	inout  nd_aib58_ch1_x0y2, 
	inout  nd_aib57_ch1_x0y2, 
	inout  nd_aib56_ch1_x0y2, 
	inout  nd_aib55_ch1_x0y2, 
	inout  nd_aib54_ch1_x0y2, 
	inout  nd_aib53_ch1_x0y2, 
	inout  nd_aib52_ch1_x0y2, 
	inout  nd_aib51_ch1_x0y2, 
	inout  nd_aib50_ch1_x0y2, 
	inout  nd_aib49_ch1_x0y2, 
	inout  nd_aib48_ch1_x0y2, 
	inout  nd_aib47_ch1_x0y2, 
	inout  nd_aib46_ch1_x0y2, 
	inout  nd_aib45_ch1_x0y2, 
	inout  nd_aib44_ch1_x0y2, 
	inout  nd_aib43_ch1_x0y2, 
	inout  nd_aib42_ch1_x0y2, 
	inout  nd_aib41_ch1_x0y2, 
	inout  nd_aib40_ch1_x0y2, 
	inout  nd_aib39_ch1_x0y2, 
	inout  nd_aib38_ch1_x0y2, 
	inout  nd_aib37_ch1_x0y2, 
	inout  nd_aib36_ch1_x0y2, 
	inout  nd_aib35_ch1_x0y2, 
	inout  nd_aib34_ch1_x0y2, 
	inout  nd_aib33_ch1_x0y2, 
	inout  nd_aib32_ch1_x0y2, 
	inout  nd_aib31_ch1_x0y2, 
	inout  nd_aib30_ch1_x0y2, 
	inout  nd_aib29_ch1_x0y2, 
	inout  nd_aib28_ch1_x0y2, 
	inout  nd_aib27_ch1_x0y2, 
	inout  nd_aib26_ch1_x0y2, 
	inout  nd_aib25_ch1_x0y2, 
	inout  nd_aib24_ch1_x0y2, 
	inout  nd_aib23_ch1_x0y2, 
	inout  nd_aib22_ch1_x0y2, 
	inout  nd_aib21_ch1_x0y2, 
	inout  nd_aib20_ch1_x0y2, 
	inout  nd_aib19_ch1_x0y2, 
	inout  nd_aib18_ch1_x0y2, 
	inout  nd_aib17_ch1_x0y2, 
	inout  nd_aib16_ch1_x0y2, 
	inout  nd_aib15_ch1_x0y2, 
	inout  nd_aib14_ch1_x0y2, 
	inout  nd_aib13_ch1_x0y2, 
	inout  nd_aib12_ch1_x0y2, 
	inout  nd_aib11_ch1_x0y2, 
	inout  nd_aib10_ch1_x0y2, 
	inout  nd_aib9_ch1_x0y2, 
	inout  nd_aib8_ch1_x0y2, 
	inout  nd_aib7_ch1_x0y2, 
	inout  nd_aib6_ch1_x0y2, 
	inout  nd_aib5_ch1_x0y2, 
	inout  nd_aib4_ch1_x0y2, 
	inout  nd_aib3_ch1_x0y2, 
	inout  nd_aib2_ch1_x0y2, 
	inout  nd_aib1_ch1_x0y2, 
	inout  nd_aib0_ch1_x0y2, 
// ## START OF ch14 ( ##
        inout [95:0] m2_ch2_aib,
 	inout  nd_aib95_ch2_x0y2, 
	inout  nd_aib94_ch2_x0y2, 
	inout  nd_aib93_ch2_x0y2, 
	inout  nd_aib92_ch2_x0y2, 
	inout  nd_aib91_ch2_x0y2, 
	inout  nd_aib90_ch2_x0y2, 
	inout  nd_aib89_ch2_x0y2, 
	inout  nd_aib88_ch2_x0y2, 
	inout  nd_aib87_ch2_x0y2, 
	inout  nd_aib86_ch2_x0y2, 
	inout  nd_aib85_ch2_x0y2, 
	inout  nd_aib84_ch2_x0y2, 
	inout  nd_aib83_ch2_x0y2, 
	inout  nd_aib82_ch2_x0y2, 
	inout  nd_aib81_ch2_x0y2, 
	inout  nd_aib80_ch2_x0y2, 
	inout  nd_aib79_ch2_x0y2, 
	inout  nd_aib78_ch2_x0y2, 
	inout  nd_aib77_ch2_x0y2, 
	inout  nd_aib76_ch2_x0y2, 
	inout  nd_aib75_ch2_x0y2, 
	inout  nd_aib74_ch2_x0y2, 
	inout  nd_aib73_ch2_x0y2, 
	inout  nd_aib72_ch2_x0y2, 
	inout  nd_aib71_ch2_x0y2, 
	inout  nd_aib70_ch2_x0y2, 
	inout  nd_aib69_ch2_x0y2, 
	inout  nd_aib68_ch2_x0y2, 
	inout  nd_aib67_ch2_x0y2, 
	inout  nd_aib66_ch2_x0y2, 
	inout  nd_aib65_ch2_x0y2, 
	inout  nd_aib64_ch2_x0y2, 
	inout  nd_aib63_ch2_x0y2, 
	inout  nd_aib62_ch2_x0y2, 
	inout  nd_aib61_ch2_x0y2, 
	inout  nd_aib60_ch2_x0y2, 
	inout  nd_aib59_ch2_x0y2, 
	inout  nd_aib58_ch2_x0y2, 
	inout  nd_aib57_ch2_x0y2, 
	inout  nd_aib56_ch2_x0y2, 
	inout  nd_aib55_ch2_x0y2, 
	inout  nd_aib54_ch2_x0y2, 
	inout  nd_aib53_ch2_x0y2, 
	inout  nd_aib52_ch2_x0y2, 
	inout  nd_aib51_ch2_x0y2, 
	inout  nd_aib50_ch2_x0y2, 
	inout  nd_aib49_ch2_x0y2, 
	inout  nd_aib48_ch2_x0y2, 
	inout  nd_aib47_ch2_x0y2, 
	inout  nd_aib46_ch2_x0y2, 
	inout  nd_aib45_ch2_x0y2, 
	inout  nd_aib44_ch2_x0y2, 
	inout  nd_aib43_ch2_x0y2, 
	inout  nd_aib42_ch2_x0y2, 
	inout  nd_aib41_ch2_x0y2, 
	inout  nd_aib40_ch2_x0y2, 
	inout  nd_aib39_ch2_x0y2, 
	inout  nd_aib38_ch2_x0y2, 
	inout  nd_aib37_ch2_x0y2, 
	inout  nd_aib36_ch2_x0y2, 
	inout  nd_aib35_ch2_x0y2, 
	inout  nd_aib34_ch2_x0y2, 
	inout  nd_aib33_ch2_x0y2, 
	inout  nd_aib32_ch2_x0y2, 
	inout  nd_aib31_ch2_x0y2, 
	inout  nd_aib30_ch2_x0y2, 
	inout  nd_aib29_ch2_x0y2, 
	inout  nd_aib28_ch2_x0y2, 
	inout  nd_aib27_ch2_x0y2, 
	inout  nd_aib26_ch2_x0y2, 
	inout  nd_aib25_ch2_x0y2, 
	inout  nd_aib24_ch2_x0y2, 
	inout  nd_aib23_ch2_x0y2, 
	inout  nd_aib22_ch2_x0y2, 
	inout  nd_aib21_ch2_x0y2, 
	inout  nd_aib20_ch2_x0y2, 
	inout  nd_aib19_ch2_x0y2, 
	inout  nd_aib18_ch2_x0y2, 
	inout  nd_aib17_ch2_x0y2, 
	inout  nd_aib16_ch2_x0y2, 
	inout  nd_aib15_ch2_x0y2, 
	inout  nd_aib14_ch2_x0y2, 
	inout  nd_aib13_ch2_x0y2, 
	inout  nd_aib12_ch2_x0y2, 
	inout  nd_aib11_ch2_x0y2, 
	inout  nd_aib10_ch2_x0y2, 
	inout  nd_aib9_ch2_x0y2, 
	inout  nd_aib8_ch2_x0y2, 
	inout  nd_aib7_ch2_x0y2, 
	inout  nd_aib6_ch2_x0y2, 
	inout  nd_aib5_ch2_x0y2, 
	inout  nd_aib4_ch2_x0y2, 
	inout  nd_aib3_ch2_x0y2, 
	inout  nd_aib2_ch2_x0y2, 
	inout  nd_aib1_ch2_x0y2, 
	inout  nd_aib0_ch2_x0y2, 
// ## START OF ch15 ( ##
        inout [95:0] m2_ch3_aib,
 	inout  nd_aib95_ch3_x0y2, 
	inout  nd_aib94_ch3_x0y2, 
	inout  nd_aib93_ch3_x0y2, 
	inout  nd_aib92_ch3_x0y2, 
	inout  nd_aib91_ch3_x0y2, 
	inout  nd_aib90_ch3_x0y2, 
	inout  nd_aib89_ch3_x0y2, 
	inout  nd_aib88_ch3_x0y2, 
	inout  nd_aib87_ch3_x0y2, 
	inout  nd_aib86_ch3_x0y2, 
	inout  nd_aib85_ch3_x0y2, 
	inout  nd_aib84_ch3_x0y2, 
	inout  nd_aib83_ch3_x0y2, 
	inout  nd_aib82_ch3_x0y2, 
	inout  nd_aib81_ch3_x0y2, 
	inout  nd_aib80_ch3_x0y2, 
	inout  nd_aib79_ch3_x0y2, 
	inout  nd_aib78_ch3_x0y2, 
	inout  nd_aib77_ch3_x0y2, 
	inout  nd_aib76_ch3_x0y2, 
	inout  nd_aib75_ch3_x0y2, 
	inout  nd_aib74_ch3_x0y2, 
	inout  nd_aib73_ch3_x0y2, 
	inout  nd_aib72_ch3_x0y2, 
	inout  nd_aib71_ch3_x0y2, 
	inout  nd_aib70_ch3_x0y2, 
	inout  nd_aib69_ch3_x0y2, 
	inout  nd_aib68_ch3_x0y2, 
	inout  nd_aib67_ch3_x0y2, 
	inout  nd_aib66_ch3_x0y2, 
	inout  nd_aib65_ch3_x0y2, 
	inout  nd_aib64_ch3_x0y2, 
	inout  nd_aib63_ch3_x0y2, 
	inout  nd_aib62_ch3_x0y2, 
	inout  nd_aib61_ch3_x0y2, 
	inout  nd_aib60_ch3_x0y2, 
	inout  nd_aib59_ch3_x0y2, 
	inout  nd_aib58_ch3_x0y2, 
	inout  nd_aib57_ch3_x0y2, 
	inout  nd_aib56_ch3_x0y2, 
	inout  nd_aib55_ch3_x0y2, 
	inout  nd_aib54_ch3_x0y2, 
	inout  nd_aib53_ch3_x0y2, 
	inout  nd_aib52_ch3_x0y2, 
	inout  nd_aib51_ch3_x0y2, 
	inout  nd_aib50_ch3_x0y2, 
	inout  nd_aib49_ch3_x0y2, 
	inout  nd_aib48_ch3_x0y2, 
	inout  nd_aib47_ch3_x0y2, 
	inout  nd_aib46_ch3_x0y2, 
	inout  nd_aib45_ch3_x0y2, 
	inout  nd_aib44_ch3_x0y2, 
	inout  nd_aib43_ch3_x0y2, 
	inout  nd_aib42_ch3_x0y2, 
	inout  nd_aib41_ch3_x0y2, 
	inout  nd_aib40_ch3_x0y2, 
	inout  nd_aib39_ch3_x0y2, 
	inout  nd_aib38_ch3_x0y2, 
	inout  nd_aib37_ch3_x0y2, 
	inout  nd_aib36_ch3_x0y2, 
	inout  nd_aib35_ch3_x0y2, 
	inout  nd_aib34_ch3_x0y2, 
	inout  nd_aib33_ch3_x0y2, 
	inout  nd_aib32_ch3_x0y2, 
	inout  nd_aib31_ch3_x0y2, 
	inout  nd_aib30_ch3_x0y2, 
	inout  nd_aib29_ch3_x0y2, 
	inout  nd_aib28_ch3_x0y2, 
	inout  nd_aib27_ch3_x0y2, 
	inout  nd_aib26_ch3_x0y2, 
	inout  nd_aib25_ch3_x0y2, 
	inout  nd_aib24_ch3_x0y2, 
	inout  nd_aib23_ch3_x0y2, 
	inout  nd_aib22_ch3_x0y2, 
	inout  nd_aib21_ch3_x0y2, 
	inout  nd_aib20_ch3_x0y2, 
	inout  nd_aib19_ch3_x0y2, 
	inout  nd_aib18_ch3_x0y2, 
	inout  nd_aib17_ch3_x0y2, 
	inout  nd_aib16_ch3_x0y2, 
	inout  nd_aib15_ch3_x0y2, 
	inout  nd_aib14_ch3_x0y2, 
	inout  nd_aib13_ch3_x0y2, 
	inout  nd_aib12_ch3_x0y2, 
	inout  nd_aib11_ch3_x0y2, 
	inout  nd_aib10_ch3_x0y2, 
	inout  nd_aib9_ch3_x0y2, 
	inout  nd_aib8_ch3_x0y2, 
	inout  nd_aib7_ch3_x0y2, 
	inout  nd_aib6_ch3_x0y2, 
	inout  nd_aib5_ch3_x0y2, 
	inout  nd_aib4_ch3_x0y2, 
	inout  nd_aib3_ch3_x0y2, 
	inout  nd_aib2_ch3_x0y2, 
	inout  nd_aib1_ch3_x0y2, 
	inout  nd_aib0_ch3_x0y2 
  );
// ## START OF  ch0 ( ##
  aliasv xaliasv95_ch0 (
    .PLUS(nd_aib95_ch0_x0y0),
    .MINUS(m0_ch0_aib[95])
   );

  aliasv xaliasv94_ch0 (
    .PLUS(nd_aib94_ch0_x0y0),
    .MINUS(m0_ch0_aib[94])
   );

  aliasv xaliasv93_ch0 (
    .PLUS(nd_aib93_ch0_x0y0),
    .MINUS(m0_ch0_aib[93])
   );

  aliasv xaliasv92_ch0 (
    .PLUS(nd_aib92_ch0_x0y0),
    .MINUS(m0_ch0_aib[92])
   );

  aliasv xaliasv91_ch0 (
    .PLUS(nd_aib91_ch0_x0y0),
    .MINUS(m0_ch0_aib[91])
   );

  aliasv xaliasv90_ch0 (
    .PLUS(nd_aib90_ch0_x0y0),
    .MINUS(m0_ch0_aib[90])
   );

  aliasv xaliasv89_ch0 (
    .PLUS(nd_aib89_ch0_x0y0),
    .MINUS(m0_ch0_aib[89])
   );

  aliasv xaliasv88_ch0 (
    .PLUS(nd_aib88_ch0_x0y0),
    .MINUS(m0_ch0_aib[88])
   );

  aliasv xaliasv87_ch0 (
    .PLUS(nd_aib87_ch0_x0y0),
    .MINUS(m0_ch0_aib[87])
   );

  aliasv xaliasv86_ch0 (
    .PLUS(nd_aib86_ch0_x0y0),
    .MINUS(m0_ch0_aib[86])
   );

  aliasv xaliasv85_ch0 (
    .PLUS(nd_aib85_ch0_x0y0),
    .MINUS(m0_ch0_aib[85])
   );

  aliasv xaliasv84_ch0 (
    .PLUS(nd_aib84_ch0_x0y0),
    .MINUS(m0_ch0_aib[84])
   );

  aliasv xaliasv83_ch0 (
    .PLUS(nd_aib83_ch0_x0y0),
    .MINUS(m0_ch0_aib[83])
   );

  aliasv xaliasv82_ch0 (
    .PLUS(nd_aib82_ch0_x0y0),
    .MINUS(m0_ch0_aib[82])
   );

  aliasv xaliasv81_ch0 (
    .PLUS(nd_aib81_ch0_x0y0),
    .MINUS(m0_ch0_aib[81])
   );

  aliasv xaliasv80_ch0 (
    .PLUS(nd_aib80_ch0_x0y0),
    .MINUS(m0_ch0_aib[80])
   );

  aliasv xaliasv79_ch0 (
    .PLUS(nd_aib79_ch0_x0y0),
    .MINUS(m0_ch0_aib[79])
   );

  aliasv xaliasv78_ch0 (
    .PLUS(nd_aib78_ch0_x0y0),
    .MINUS(m0_ch0_aib[78])
   );

  aliasv xaliasv77_ch0 (
    .PLUS(nd_aib77_ch0_x0y0),
    .MINUS(m0_ch0_aib[77])
   );

  aliasv xaliasv76_ch0 (
    .PLUS(nd_aib76_ch0_x0y0),
    .MINUS(m0_ch0_aib[76])
   );

  aliasv xaliasv75_ch0 (
    .PLUS(nd_aib75_ch0_x0y0),
    .MINUS(m0_ch0_aib[75])
   );

  aliasv xaliasv74_ch0 (
    .PLUS(nd_aib74_ch0_x0y0),
    .MINUS(m0_ch0_aib[74])
   );

  aliasv xaliasv73_ch0 (
    .PLUS(nd_aib73_ch0_x0y0),
    .MINUS(m0_ch0_aib[73])
   );

  aliasv xaliasv72_ch0 (
    .PLUS(nd_aib72_ch0_x0y0),
    .MINUS(m0_ch0_aib[72])
   );

  aliasv xaliasv71_ch0 (
    .PLUS(nd_aib71_ch0_x0y0),
    .MINUS(m0_ch0_aib[71])
   );

  aliasv xaliasv70_ch0 (
    .PLUS(nd_aib70_ch0_x0y0),
    .MINUS(m0_ch0_aib[70])
   );

  aliasv xaliasv69_ch0 (
    .PLUS(nd_aib69_ch0_x0y0),
    .MINUS(m0_ch0_aib[69])
   );

  aliasv xaliasv68_ch0 (
    .PLUS(nd_aib68_ch0_x0y0),
    .MINUS(m0_ch0_aib[68])
   );

  aliasv xaliasv67_ch0 (
    .PLUS(nd_aib67_ch0_x0y0),
    .MINUS(m0_ch0_aib[67])
   );

  aliasv xaliasv66_ch0 (
    .PLUS(nd_aib66_ch0_x0y0),
    .MINUS(m0_ch0_aib[66])
   );

  aliasv xaliasv65_ch0 (
    .PLUS(nd_aib65_ch0_x0y0),
    .MINUS(m0_ch0_aib[65])
   );

  aliasv xaliasv64_ch0 (
    .PLUS(nd_aib64_ch0_x0y0),
    .MINUS(m0_ch0_aib[64])
   );

  aliasv xaliasv63_ch0 (
    .PLUS(nd_aib63_ch0_x0y0),
    .MINUS(m0_ch0_aib[63])
   );

  aliasv xaliasv62_ch0 (
    .PLUS(nd_aib62_ch0_x0y0),
    .MINUS(m0_ch0_aib[62])
   );

  aliasv xaliasv61_ch0 (
    .PLUS(nd_aib61_ch0_x0y0),
    .MINUS(m0_ch0_aib[61])
   );

  aliasv xaliasv60_ch0 (
    .PLUS(nd_aib60_ch0_x0y0),
    .MINUS(m0_ch0_aib[60])
   );

  aliasv xaliasv59_ch0 (
    .PLUS(nd_aib59_ch0_x0y0),
    .MINUS(m0_ch0_aib[59])
   );

  aliasv xaliasv58_ch0 (
    .PLUS(nd_aib58_ch0_x0y0),
    .MINUS(m0_ch0_aib[58])
   );

  aliasv xaliasv57_ch0 (
    .PLUS(nd_aib57_ch0_x0y0),
    .MINUS(m0_ch0_aib[57])
   );

  aliasv xaliasv56_ch0 (
    .PLUS(nd_aib56_ch0_x0y0),
    .MINUS(m0_ch0_aib[56])
   );

  aliasv xaliasv55_ch0 (
    .PLUS(nd_aib55_ch0_x0y0),
    .MINUS(m0_ch0_aib[55])
   );

  aliasv xaliasv54_ch0 (
    .PLUS(nd_aib54_ch0_x0y0),
    .MINUS(m0_ch0_aib[54])
   );

  aliasv xaliasv53_ch0 (
    .PLUS(nd_aib53_ch0_x0y0),
    .MINUS(m0_ch0_aib[53])
   );

  aliasv xaliasv52_ch0 (
    .PLUS(nd_aib52_ch0_x0y0),
    .MINUS(m0_ch0_aib[52])
   );

  aliasv xaliasv51_ch0 (
    .PLUS(nd_aib51_ch0_x0y0),
    .MINUS(m0_ch0_aib[51])
   );

  aliasv xaliasv50_ch0 (
    .PLUS(nd_aib50_ch0_x0y0),
    .MINUS(m0_ch0_aib[50])
   );

  aliasv xaliasv49_ch0 (
    .PLUS(nd_aib49_ch0_x0y0),
    .MINUS(m0_ch0_aib[49])
   );

  aliasv xaliasv48_ch0 (
    .PLUS(nd_aib48_ch0_x0y0),
    .MINUS(m0_ch0_aib[48])
   );

  aliasv xaliasv47_ch0 (
    .PLUS(nd_aib47_ch0_x0y0),
    .MINUS(m0_ch0_aib[47])
   );

  aliasv xaliasv46_ch0 (
    .PLUS(nd_aib46_ch0_x0y0),
    .MINUS(m0_ch0_aib[46])
   );

  aliasv xaliasv45_ch0 (
    .PLUS(nd_aib45_ch0_x0y0),
    .MINUS(m0_ch0_aib[45])
   );

  aliasv xaliasv44_ch0 (
    .PLUS(nd_aib44_ch0_x0y0),
    .MINUS(m0_ch0_aib[44])
   );

  aliasv xaliasv43_ch0 (
    .PLUS(nd_aib43_ch0_x0y0),
    .MINUS(m0_ch0_aib[43])
   );

  aliasv xaliasv42_ch0 (
    .PLUS(nd_aib42_ch0_x0y0),
    .MINUS(m0_ch0_aib[42])
   );

  aliasv xaliasv41_ch0 (
    .PLUS(nd_aib41_ch0_x0y0),
    .MINUS(m0_ch0_aib[41])
   );

  aliasv xaliasv40_ch0 (
    .PLUS(nd_aib40_ch0_x0y0),
    .MINUS(m0_ch0_aib[40])
   );

  aliasv xaliasv39_ch0 (
    .PLUS(nd_aib39_ch0_x0y0),
    .MINUS(m0_ch0_aib[39])
   );

  aliasv xaliasv38_ch0 (
    .PLUS(nd_aib38_ch0_x0y0),
    .MINUS(m0_ch0_aib[38])
   );

  aliasv xaliasv37_ch0 (
    .PLUS(nd_aib37_ch0_x0y0),
    .MINUS(m0_ch0_aib[37])
   );

  aliasv xaliasv36_ch0 (
    .PLUS(nd_aib36_ch0_x0y0),
    .MINUS(m0_ch0_aib[36])
   );

  aliasv xaliasv35_ch0 (
    .PLUS(nd_aib35_ch0_x0y0),
    .MINUS(m0_ch0_aib[35])
   );

  aliasv xaliasv34_ch0 (
    .PLUS(nd_aib34_ch0_x0y0),
    .MINUS(m0_ch0_aib[34])
   );

  aliasv xaliasv33_ch0 (
    .PLUS(nd_aib33_ch0_x0y0),
    .MINUS(m0_ch0_aib[33])
   );

  aliasv xaliasv32_ch0 (
    .PLUS(nd_aib32_ch0_x0y0),
    .MINUS(m0_ch0_aib[32])
   );

  aliasv xaliasv31_ch0 (
    .PLUS(nd_aib31_ch0_x0y0),
    .MINUS(m0_ch0_aib[31])
   );

  aliasv xaliasv30_ch0 (
    .PLUS(nd_aib30_ch0_x0y0),
    .MINUS(m0_ch0_aib[30])
   );

  aliasv xaliasv29_ch0 (
    .PLUS(nd_aib29_ch0_x0y0),
    .MINUS(m0_ch0_aib[29])
   );

  aliasv xaliasv28_ch0 (
    .PLUS(nd_aib28_ch0_x0y0),
    .MINUS(m0_ch0_aib[28])
   );

  aliasv xaliasv27_ch0 (
    .PLUS(nd_aib27_ch0_x0y0),
    .MINUS(m0_ch0_aib[27])
   );

  aliasv xaliasv26_ch0 (
    .PLUS(nd_aib26_ch0_x0y0),
    .MINUS(m0_ch0_aib[26])
   );

  aliasv xaliasv25_ch0 (
    .PLUS(nd_aib25_ch0_x0y0),
    .MINUS(m0_ch0_aib[25])
   );

  aliasv xaliasv24_ch0 (
    .PLUS(nd_aib24_ch0_x0y0),
    .MINUS(m0_ch0_aib[24])
   );

  aliasv xaliasv23_ch0 (
    .PLUS(nd_aib23_ch0_x0y0),
    .MINUS(m0_ch0_aib[23])
   );

  aliasv xaliasv22_ch0 (
    .PLUS(nd_aib22_ch0_x0y0),
    .MINUS(m0_ch0_aib[22])
   );

  aliasv xaliasv21_ch0 (
    .PLUS(nd_aib21_ch0_x0y0),
    .MINUS(m0_ch0_aib[21])
   );

  aliasv xaliasv20_ch0 (
    .PLUS(nd_aib20_ch0_x0y0),
    .MINUS(m0_ch0_aib[20])
   );

  aliasv xaliasv19_ch0 (
    .PLUS(nd_aib19_ch0_x0y0),
    .MINUS(m0_ch0_aib[19])
   );

  aliasv xaliasv18_ch0 (
    .PLUS(nd_aib18_ch0_x0y0),
    .MINUS(m0_ch0_aib[18])
   );

  aliasv xaliasv17_ch0 (
    .PLUS(nd_aib17_ch0_x0y0),
    .MINUS(m0_ch0_aib[17])
   );

  aliasv xaliasv16_ch0 (
    .PLUS(nd_aib16_ch0_x0y0),
    .MINUS(m0_ch0_aib[16])
   );

  aliasv xaliasv15_ch0 (
    .PLUS(nd_aib15_ch0_x0y0),
    .MINUS(m0_ch0_aib[15])
   );

  aliasv xaliasv14_ch0 (
    .PLUS(nd_aib14_ch0_x0y0),
    .MINUS(m0_ch0_aib[14])
   );

  aliasv xaliasv13_ch0 (
    .PLUS(nd_aib13_ch0_x0y0),
    .MINUS(m0_ch0_aib[13])
   );

  aliasv xaliasv12_ch0 (
    .PLUS(nd_aib12_ch0_x0y0),
    .MINUS(m0_ch0_aib[12])
   );

  aliasv xaliasv11_ch0 (
    .PLUS(nd_aib11_ch0_x0y0),
    .MINUS(m0_ch0_aib[11])
   );

  aliasv xaliasv10_ch0 (
    .PLUS(nd_aib10_ch0_x0y0),
    .MINUS(m0_ch0_aib[10])
   );

  aliasv xaliasv9_ch0 (
    .PLUS(nd_aib9_ch0_x0y0),
    .MINUS(m0_ch0_aib[9])
   );

  aliasv xaliasv8_ch0 (
    .PLUS(nd_aib8_ch0_x0y0),
    .MINUS(m0_ch0_aib[8])
   );

  aliasv xaliasv7_ch0 (
    .PLUS(nd_aib7_ch0_x0y0),
    .MINUS(m0_ch0_aib[7])
   );

  aliasv xaliasv6_ch0 (
    .PLUS(nd_aib6_ch0_x0y0),
    .MINUS(m0_ch0_aib[6])
   );

  aliasv xaliasv5_ch0 (
    .PLUS(nd_aib5_ch0_x0y0),
    .MINUS(m0_ch0_aib[5])
   );

  aliasv xaliasv4_ch0 (
    .PLUS(nd_aib4_ch0_x0y0),
    .MINUS(m0_ch0_aib[4])
   );

  aliasv xaliasv3_ch0 (
    .PLUS(nd_aib3_ch0_x0y0),
    .MINUS(m0_ch0_aib[3])
   );

  aliasv xaliasv2_ch0 (
    .PLUS(nd_aib2_ch0_x0y0),
    .MINUS(m0_ch0_aib[2])
   );

  aliasv xaliasv1_ch0 (
    .PLUS(nd_aib1_ch0_x0y0),
    .MINUS(m0_ch0_aib[1])
   );

  aliasv xaliasv0_ch0 (
    .PLUS(nd_aib0_ch0_x0y0),
    .MINUS(m0_ch0_aib[0])
   );

// ## START OF  ch1 ( ##
  aliasv xaliasv95_ch1 (
    .PLUS(nd_aib95_ch1_x0y0),
    .MINUS(m0_ch1_aib[95])
   );

  aliasv xaliasv94_ch1 (
    .PLUS(nd_aib94_ch1_x0y0),
    .MINUS(m0_ch1_aib[94])
   );

  aliasv xaliasv93_ch1 (
    .PLUS(nd_aib93_ch1_x0y0),
    .MINUS(m0_ch1_aib[93])
   );

  aliasv xaliasv92_ch1 (
    .PLUS(nd_aib92_ch1_x0y0),
    .MINUS(m0_ch1_aib[92])
   );

  aliasv xaliasv91_ch1 (
    .PLUS(nd_aib91_ch1_x0y0),
    .MINUS(m0_ch1_aib[91])
   );

  aliasv xaliasv90_ch1 (
    .PLUS(nd_aib90_ch1_x0y0),
    .MINUS(m0_ch1_aib[90])
   );

  aliasv xaliasv89_ch1 (
    .PLUS(nd_aib89_ch1_x0y0),
    .MINUS(m0_ch1_aib[89])
   );

  aliasv xaliasv88_ch1 (
    .PLUS(nd_aib88_ch1_x0y0),
    .MINUS(m0_ch1_aib[88])
   );

  aliasv xaliasv87_ch1 (
    .PLUS(nd_aib87_ch1_x0y0),
    .MINUS(m0_ch1_aib[87])
   );

  aliasv xaliasv86_ch1 (
    .PLUS(nd_aib86_ch1_x0y0),
    .MINUS(m0_ch1_aib[86])
   );

  aliasv xaliasv85_ch1 (
    .PLUS(nd_aib85_ch1_x0y0),
    .MINUS(m0_ch1_aib[85])
   );

  aliasv xaliasv84_ch1 (
    .PLUS(nd_aib84_ch1_x0y0),
    .MINUS(m0_ch1_aib[84])
   );

  aliasv xaliasv83_ch1 (
    .PLUS(nd_aib83_ch1_x0y0),
    .MINUS(m0_ch1_aib[83])
   );

  aliasv xaliasv82_ch1 (
    .PLUS(nd_aib82_ch1_x0y0),
    .MINUS(m0_ch1_aib[82])
   );

  aliasv xaliasv81_ch1 (
    .PLUS(nd_aib81_ch1_x0y0),
    .MINUS(m0_ch1_aib[81])
   );

  aliasv xaliasv80_ch1 (
    .PLUS(nd_aib80_ch1_x0y0),
    .MINUS(m0_ch1_aib[80])
   );

  aliasv xaliasv79_ch1 (
    .PLUS(nd_aib79_ch1_x0y0),
    .MINUS(m0_ch1_aib[79])
   );

  aliasv xaliasv78_ch1 (
    .PLUS(nd_aib78_ch1_x0y0),
    .MINUS(m0_ch1_aib[78])
   );

  aliasv xaliasv77_ch1 (
    .PLUS(nd_aib77_ch1_x0y0),
    .MINUS(m0_ch1_aib[77])
   );

  aliasv xaliasv76_ch1 (
    .PLUS(nd_aib76_ch1_x0y0),
    .MINUS(m0_ch1_aib[76])
   );

  aliasv xaliasv75_ch1 (
    .PLUS(nd_aib75_ch1_x0y0),
    .MINUS(m0_ch1_aib[75])
   );

  aliasv xaliasv74_ch1 (
    .PLUS(nd_aib74_ch1_x0y0),
    .MINUS(m0_ch1_aib[74])
   );

  aliasv xaliasv73_ch1 (
    .PLUS(nd_aib73_ch1_x0y0),
    .MINUS(m0_ch1_aib[73])
   );

  aliasv xaliasv72_ch1 (
    .PLUS(nd_aib72_ch1_x0y0),
    .MINUS(m0_ch1_aib[72])
   );

  aliasv xaliasv71_ch1 (
    .PLUS(nd_aib71_ch1_x0y0),
    .MINUS(m0_ch1_aib[71])
   );

  aliasv xaliasv70_ch1 (
    .PLUS(nd_aib70_ch1_x0y0),
    .MINUS(m0_ch1_aib[70])
   );

  aliasv xaliasv69_ch1 (
    .PLUS(nd_aib69_ch1_x0y0),
    .MINUS(m0_ch1_aib[69])
   );

  aliasv xaliasv68_ch1 (
    .PLUS(nd_aib68_ch1_x0y0),
    .MINUS(m0_ch1_aib[68])
   );

  aliasv xaliasv67_ch1 (
    .PLUS(nd_aib67_ch1_x0y0),
    .MINUS(m0_ch1_aib[67])
   );

  aliasv xaliasv66_ch1 (
    .PLUS(nd_aib66_ch1_x0y0),
    .MINUS(m0_ch1_aib[66])
   );

  aliasv xaliasv65_ch1 (
    .PLUS(nd_aib65_ch1_x0y0),
    .MINUS(m0_ch1_aib[65])
   );

  aliasv xaliasv64_ch1 (
    .PLUS(nd_aib64_ch1_x0y0),
    .MINUS(m0_ch1_aib[64])
   );

  aliasv xaliasv63_ch1 (
    .PLUS(nd_aib63_ch1_x0y0),
    .MINUS(m0_ch1_aib[63])
   );

  aliasv xaliasv62_ch1 (
    .PLUS(nd_aib62_ch1_x0y0),
    .MINUS(m0_ch1_aib[62])
   );

  aliasv xaliasv61_ch1 (
    .PLUS(nd_aib61_ch1_x0y0),
    .MINUS(m0_ch1_aib[61])
   );

  aliasv xaliasv60_ch1 (
    .PLUS(nd_aib60_ch1_x0y0),
    .MINUS(m0_ch1_aib[60])
   );

  aliasv xaliasv59_ch1 (
    .PLUS(nd_aib59_ch1_x0y0),
    .MINUS(m0_ch1_aib[59])
   );

  aliasv xaliasv58_ch1 (
    .PLUS(nd_aib58_ch1_x0y0),
    .MINUS(m0_ch1_aib[58])
   );

  aliasv xaliasv57_ch1 (
    .PLUS(nd_aib57_ch1_x0y0),
    .MINUS(m0_ch1_aib[57])
   );

  aliasv xaliasv56_ch1 (
    .PLUS(nd_aib56_ch1_x0y0),
    .MINUS(m0_ch1_aib[56])
   );

  aliasv xaliasv55_ch1 (
    .PLUS(nd_aib55_ch1_x0y0),
    .MINUS(m0_ch1_aib[55])
   );

  aliasv xaliasv54_ch1 (
    .PLUS(nd_aib54_ch1_x0y0),
    .MINUS(m0_ch1_aib[54])
   );

  aliasv xaliasv53_ch1 (
    .PLUS(nd_aib53_ch1_x0y0),
    .MINUS(m0_ch1_aib[53])
   );

  aliasv xaliasv52_ch1 (
    .PLUS(nd_aib52_ch1_x0y0),
    .MINUS(m0_ch1_aib[52])
   );

  aliasv xaliasv51_ch1 (
    .PLUS(nd_aib51_ch1_x0y0),
    .MINUS(m0_ch1_aib[51])
   );

  aliasv xaliasv50_ch1 (
    .PLUS(nd_aib50_ch1_x0y0),
    .MINUS(m0_ch1_aib[50])
   );

  aliasv xaliasv49_ch1 (
    .PLUS(nd_aib49_ch1_x0y0),
    .MINUS(m0_ch1_aib[49])
   );

  aliasv xaliasv48_ch1 (
    .PLUS(nd_aib48_ch1_x0y0),
    .MINUS(m0_ch1_aib[48])
   );

  aliasv xaliasv47_ch1 (
    .PLUS(nd_aib47_ch1_x0y0),
    .MINUS(m0_ch1_aib[47])
   );

  aliasv xaliasv46_ch1 (
    .PLUS(nd_aib46_ch1_x0y0),
    .MINUS(m0_ch1_aib[46])
   );

  aliasv xaliasv45_ch1 (
    .PLUS(nd_aib45_ch1_x0y0),
    .MINUS(m0_ch1_aib[45])
   );

  aliasv xaliasv44_ch1 (
    .PLUS(nd_aib44_ch1_x0y0),
    .MINUS(m0_ch1_aib[44])
   );

  aliasv xaliasv43_ch1 (
    .PLUS(nd_aib43_ch1_x0y0),
    .MINUS(m0_ch1_aib[43])
   );

  aliasv xaliasv42_ch1 (
    .PLUS(nd_aib42_ch1_x0y0),
    .MINUS(m0_ch1_aib[42])
   );

  aliasv xaliasv41_ch1 (
    .PLUS(nd_aib41_ch1_x0y0),
    .MINUS(m0_ch1_aib[41])
   );

  aliasv xaliasv40_ch1 (
    .PLUS(nd_aib40_ch1_x0y0),
    .MINUS(m0_ch1_aib[40])
   );

  aliasv xaliasv39_ch1 (
    .PLUS(nd_aib39_ch1_x0y0),
    .MINUS(m0_ch1_aib[39])
   );

  aliasv xaliasv38_ch1 (
    .PLUS(nd_aib38_ch1_x0y0),
    .MINUS(m0_ch1_aib[38])
   );

  aliasv xaliasv37_ch1 (
    .PLUS(nd_aib37_ch1_x0y0),
    .MINUS(m0_ch1_aib[37])
   );

  aliasv xaliasv36_ch1 (
    .PLUS(nd_aib36_ch1_x0y0),
    .MINUS(m0_ch1_aib[36])
   );

  aliasv xaliasv35_ch1 (
    .PLUS(nd_aib35_ch1_x0y0),
    .MINUS(m0_ch1_aib[35])
   );

  aliasv xaliasv34_ch1 (
    .PLUS(nd_aib34_ch1_x0y0),
    .MINUS(m0_ch1_aib[34])
   );

  aliasv xaliasv33_ch1 (
    .PLUS(nd_aib33_ch1_x0y0),
    .MINUS(m0_ch1_aib[33])
   );

  aliasv xaliasv32_ch1 (
    .PLUS(nd_aib32_ch1_x0y0),
    .MINUS(m0_ch1_aib[32])
   );

  aliasv xaliasv31_ch1 (
    .PLUS(nd_aib31_ch1_x0y0),
    .MINUS(m0_ch1_aib[31])
   );

  aliasv xaliasv30_ch1 (
    .PLUS(nd_aib30_ch1_x0y0),
    .MINUS(m0_ch1_aib[30])
   );

  aliasv xaliasv29_ch1 (
    .PLUS(nd_aib29_ch1_x0y0),
    .MINUS(m0_ch1_aib[29])
   );

  aliasv xaliasv28_ch1 (
    .PLUS(nd_aib28_ch1_x0y0),
    .MINUS(m0_ch1_aib[28])
   );

  aliasv xaliasv27_ch1 (
    .PLUS(nd_aib27_ch1_x0y0),
    .MINUS(m0_ch1_aib[27])
   );

  aliasv xaliasv26_ch1 (
    .PLUS(nd_aib26_ch1_x0y0),
    .MINUS(m0_ch1_aib[26])
   );

  aliasv xaliasv25_ch1 (
    .PLUS(nd_aib25_ch1_x0y0),
    .MINUS(m0_ch1_aib[25])
   );

  aliasv xaliasv24_ch1 (
    .PLUS(nd_aib24_ch1_x0y0),
    .MINUS(m0_ch1_aib[24])
   );

  aliasv xaliasv23_ch1 (
    .PLUS(nd_aib23_ch1_x0y0),
    .MINUS(m0_ch1_aib[23])
   );

  aliasv xaliasv22_ch1 (
    .PLUS(nd_aib22_ch1_x0y0),
    .MINUS(m0_ch1_aib[22])
   );

  aliasv xaliasv21_ch1 (
    .PLUS(nd_aib21_ch1_x0y0),
    .MINUS(m0_ch1_aib[21])
   );

  aliasv xaliasv20_ch1 (
    .PLUS(nd_aib20_ch1_x0y0),
    .MINUS(m0_ch1_aib[20])
   );

  aliasv xaliasv19_ch1 (
    .PLUS(nd_aib19_ch1_x0y0),
    .MINUS(m0_ch1_aib[19])
   );

  aliasv xaliasv18_ch1 (
    .PLUS(nd_aib18_ch1_x0y0),
    .MINUS(m0_ch1_aib[18])
   );

  aliasv xaliasv17_ch1 (
    .PLUS(nd_aib17_ch1_x0y0),
    .MINUS(m0_ch1_aib[17])
   );

  aliasv xaliasv16_ch1 (
    .PLUS(nd_aib16_ch1_x0y0),
    .MINUS(m0_ch1_aib[16])
   );

  aliasv xaliasv15_ch1 (
    .PLUS(nd_aib15_ch1_x0y0),
    .MINUS(m0_ch1_aib[15])
   );

  aliasv xaliasv14_ch1 (
    .PLUS(nd_aib14_ch1_x0y0),
    .MINUS(m0_ch1_aib[14])
   );

  aliasv xaliasv13_ch1 (
    .PLUS(nd_aib13_ch1_x0y0),
    .MINUS(m0_ch1_aib[13])
   );

  aliasv xaliasv12_ch1 (
    .PLUS(nd_aib12_ch1_x0y0),
    .MINUS(m0_ch1_aib[12])
   );

  aliasv xaliasv11_ch1 (
    .PLUS(nd_aib11_ch1_x0y0),
    .MINUS(m0_ch1_aib[11])
   );

  aliasv xaliasv10_ch1 (
    .PLUS(nd_aib10_ch1_x0y0),
    .MINUS(m0_ch1_aib[10])
   );

  aliasv xaliasv9_ch1 (
    .PLUS(nd_aib9_ch1_x0y0),
    .MINUS(m0_ch1_aib[9])
   );

  aliasv xaliasv8_ch1 (
    .PLUS(nd_aib8_ch1_x0y0),
    .MINUS(m0_ch1_aib[8])
   );

  aliasv xaliasv7_ch1 (
    .PLUS(nd_aib7_ch1_x0y0),
    .MINUS(m0_ch1_aib[7])
   );

  aliasv xaliasv6_ch1 (
    .PLUS(nd_aib6_ch1_x0y0),
    .MINUS(m0_ch1_aib[6])
   );

  aliasv xaliasv5_ch1 (
    .PLUS(nd_aib5_ch1_x0y0),
    .MINUS(m0_ch1_aib[5])
   );

  aliasv xaliasv4_ch1 (
    .PLUS(nd_aib4_ch1_x0y0),
    .MINUS(m0_ch1_aib[4])
   );

  aliasv xaliasv3_ch1 (
    .PLUS(nd_aib3_ch1_x0y0),
    .MINUS(m0_ch1_aib[3])
   );

  aliasv xaliasv2_ch1 (
    .PLUS(nd_aib2_ch1_x0y0),
    .MINUS(m0_ch1_aib[2])
   );

  aliasv xaliasv1_ch1 (
    .PLUS(nd_aib1_ch1_x0y0),
    .MINUS(m0_ch1_aib[1])
   );

  aliasv xaliasv0_ch1 (
    .PLUS(nd_aib0_ch1_x0y0),
    .MINUS(m0_ch1_aib[0])
   );

// ## START OF  ch2 ( ##
  aliasv xaliasv95_ch2 (
    .PLUS(nd_aib95_ch2_x0y0),
    .MINUS(m0_ch2_aib[95])
   );

  aliasv xaliasv94_ch2 (
    .PLUS(nd_aib94_ch2_x0y0),
    .MINUS(m0_ch2_aib[94])
   );

  aliasv xaliasv93_ch2 (
    .PLUS(nd_aib93_ch2_x0y0),
    .MINUS(m0_ch2_aib[93])
   );

  aliasv xaliasv92_ch2 (
    .PLUS(nd_aib92_ch2_x0y0),
    .MINUS(m0_ch2_aib[92])
   );

  aliasv xaliasv91_ch2 (
    .PLUS(nd_aib91_ch2_x0y0),
    .MINUS(m0_ch2_aib[91])
   );

  aliasv xaliasv90_ch2 (
    .PLUS(nd_aib90_ch2_x0y0),
    .MINUS(m0_ch2_aib[90])
   );

  aliasv xaliasv89_ch2 (
    .PLUS(nd_aib89_ch2_x0y0),
    .MINUS(m0_ch2_aib[89])
   );

  aliasv xaliasv88_ch2 (
    .PLUS(nd_aib88_ch2_x0y0),
    .MINUS(m0_ch2_aib[88])
   );

  aliasv xaliasv87_ch2 (
    .PLUS(nd_aib87_ch2_x0y0),
    .MINUS(m0_ch2_aib[87])
   );

  aliasv xaliasv86_ch2 (
    .PLUS(nd_aib86_ch2_x0y0),
    .MINUS(m0_ch2_aib[86])
   );

  aliasv xaliasv85_ch2 (
    .PLUS(nd_aib85_ch2_x0y0),
    .MINUS(m0_ch2_aib[85])
   );

  aliasv xaliasv84_ch2 (
    .PLUS(nd_aib84_ch2_x0y0),
    .MINUS(m0_ch2_aib[84])
   );

  aliasv xaliasv83_ch2 (
    .PLUS(nd_aib83_ch2_x0y0),
    .MINUS(m0_ch2_aib[83])
   );

  aliasv xaliasv82_ch2 (
    .PLUS(nd_aib82_ch2_x0y0),
    .MINUS(m0_ch2_aib[82])
   );

  aliasv xaliasv81_ch2 (
    .PLUS(nd_aib81_ch2_x0y0),
    .MINUS(m0_ch2_aib[81])
   );

  aliasv xaliasv80_ch2 (
    .PLUS(nd_aib80_ch2_x0y0),
    .MINUS(m0_ch2_aib[80])
   );

  aliasv xaliasv79_ch2 (
    .PLUS(nd_aib79_ch2_x0y0),
    .MINUS(m0_ch2_aib[79])
   );

  aliasv xaliasv78_ch2 (
    .PLUS(nd_aib78_ch2_x0y0),
    .MINUS(m0_ch2_aib[78])
   );

  aliasv xaliasv77_ch2 (
    .PLUS(nd_aib77_ch2_x0y0),
    .MINUS(m0_ch2_aib[77])
   );

  aliasv xaliasv76_ch2 (
    .PLUS(nd_aib76_ch2_x0y0),
    .MINUS(m0_ch2_aib[76])
   );

  aliasv xaliasv75_ch2 (
    .PLUS(nd_aib75_ch2_x0y0),
    .MINUS(m0_ch2_aib[75])
   );

  aliasv xaliasv74_ch2 (
    .PLUS(nd_aib74_ch2_x0y0),
    .MINUS(m0_ch2_aib[74])
   );

  aliasv xaliasv73_ch2 (
    .PLUS(nd_aib73_ch2_x0y0),
    .MINUS(m0_ch2_aib[73])
   );

  aliasv xaliasv72_ch2 (
    .PLUS(nd_aib72_ch2_x0y0),
    .MINUS(m0_ch2_aib[72])
   );

  aliasv xaliasv71_ch2 (
    .PLUS(nd_aib71_ch2_x0y0),
    .MINUS(m0_ch2_aib[71])
   );

  aliasv xaliasv70_ch2 (
    .PLUS(nd_aib70_ch2_x0y0),
    .MINUS(m0_ch2_aib[70])
   );

  aliasv xaliasv69_ch2 (
    .PLUS(nd_aib69_ch2_x0y0),
    .MINUS(m0_ch2_aib[69])
   );

  aliasv xaliasv68_ch2 (
    .PLUS(nd_aib68_ch2_x0y0),
    .MINUS(m0_ch2_aib[68])
   );

  aliasv xaliasv67_ch2 (
    .PLUS(nd_aib67_ch2_x0y0),
    .MINUS(m0_ch2_aib[67])
   );

  aliasv xaliasv66_ch2 (
    .PLUS(nd_aib66_ch2_x0y0),
    .MINUS(m0_ch2_aib[66])
   );

  aliasv xaliasv65_ch2 (
    .PLUS(nd_aib65_ch2_x0y0),
    .MINUS(m0_ch2_aib[65])
   );

  aliasv xaliasv64_ch2 (
    .PLUS(nd_aib64_ch2_x0y0),
    .MINUS(m0_ch2_aib[64])
   );

  aliasv xaliasv63_ch2 (
    .PLUS(nd_aib63_ch2_x0y0),
    .MINUS(m0_ch2_aib[63])
   );

  aliasv xaliasv62_ch2 (
    .PLUS(nd_aib62_ch2_x0y0),
    .MINUS(m0_ch2_aib[62])
   );

  aliasv xaliasv61_ch2 (
    .PLUS(nd_aib61_ch2_x0y0),
    .MINUS(m0_ch2_aib[61])
   );

  aliasv xaliasv60_ch2 (
    .PLUS(nd_aib60_ch2_x0y0),
    .MINUS(m0_ch2_aib[60])
   );

  aliasv xaliasv59_ch2 (
    .PLUS(nd_aib59_ch2_x0y0),
    .MINUS(m0_ch2_aib[59])
   );

  aliasv xaliasv58_ch2 (
    .PLUS(nd_aib58_ch2_x0y0),
    .MINUS(m0_ch2_aib[58])
   );

  aliasv xaliasv57_ch2 (
    .PLUS(nd_aib57_ch2_x0y0),
    .MINUS(m0_ch2_aib[57])
   );

  aliasv xaliasv56_ch2 (
    .PLUS(nd_aib56_ch2_x0y0),
    .MINUS(m0_ch2_aib[56])
   );

  aliasv xaliasv55_ch2 (
    .PLUS(nd_aib55_ch2_x0y0),
    .MINUS(m0_ch2_aib[55])
   );

  aliasv xaliasv54_ch2 (
    .PLUS(nd_aib54_ch2_x0y0),
    .MINUS(m0_ch2_aib[54])
   );

  aliasv xaliasv53_ch2 (
    .PLUS(nd_aib53_ch2_x0y0),
    .MINUS(m0_ch2_aib[53])
   );

  aliasv xaliasv52_ch2 (
    .PLUS(nd_aib52_ch2_x0y0),
    .MINUS(m0_ch2_aib[52])
   );

  aliasv xaliasv51_ch2 (
    .PLUS(nd_aib51_ch2_x0y0),
    .MINUS(m0_ch2_aib[51])
   );

  aliasv xaliasv50_ch2 (
    .PLUS(nd_aib50_ch2_x0y0),
    .MINUS(m0_ch2_aib[50])
   );

  aliasv xaliasv49_ch2 (
    .PLUS(nd_aib49_ch2_x0y0),
    .MINUS(m0_ch2_aib[49])
   );

  aliasv xaliasv48_ch2 (
    .PLUS(nd_aib48_ch2_x0y0),
    .MINUS(m0_ch2_aib[48])
   );

  aliasv xaliasv47_ch2 (
    .PLUS(nd_aib47_ch2_x0y0),
    .MINUS(m0_ch2_aib[47])
   );

  aliasv xaliasv46_ch2 (
    .PLUS(nd_aib46_ch2_x0y0),
    .MINUS(m0_ch2_aib[46])
   );

  aliasv xaliasv45_ch2 (
    .PLUS(nd_aib45_ch2_x0y0),
    .MINUS(m0_ch2_aib[45])
   );

  aliasv xaliasv44_ch2 (
    .PLUS(nd_aib44_ch2_x0y0),
    .MINUS(m0_ch2_aib[44])
   );

  aliasv xaliasv43_ch2 (
    .PLUS(nd_aib43_ch2_x0y0),
    .MINUS(m0_ch2_aib[43])
   );

  aliasv xaliasv42_ch2 (
    .PLUS(nd_aib42_ch2_x0y0),
    .MINUS(m0_ch2_aib[42])
   );

  aliasv xaliasv41_ch2 (
    .PLUS(nd_aib41_ch2_x0y0),
    .MINUS(m0_ch2_aib[41])
   );

  aliasv xaliasv40_ch2 (
    .PLUS(nd_aib40_ch2_x0y0),
    .MINUS(m0_ch2_aib[40])
   );

  aliasv xaliasv39_ch2 (
    .PLUS(nd_aib39_ch2_x0y0),
    .MINUS(m0_ch2_aib[39])
   );

  aliasv xaliasv38_ch2 (
    .PLUS(nd_aib38_ch2_x0y0),
    .MINUS(m0_ch2_aib[38])
   );

  aliasv xaliasv37_ch2 (
    .PLUS(nd_aib37_ch2_x0y0),
    .MINUS(m0_ch2_aib[37])
   );

  aliasv xaliasv36_ch2 (
    .PLUS(nd_aib36_ch2_x0y0),
    .MINUS(m0_ch2_aib[36])
   );

  aliasv xaliasv35_ch2 (
    .PLUS(nd_aib35_ch2_x0y0),
    .MINUS(m0_ch2_aib[35])
   );

  aliasv xaliasv34_ch2 (
    .PLUS(nd_aib34_ch2_x0y0),
    .MINUS(m0_ch2_aib[34])
   );

  aliasv xaliasv33_ch2 (
    .PLUS(nd_aib33_ch2_x0y0),
    .MINUS(m0_ch2_aib[33])
   );

  aliasv xaliasv32_ch2 (
    .PLUS(nd_aib32_ch2_x0y0),
    .MINUS(m0_ch2_aib[32])
   );

  aliasv xaliasv31_ch2 (
    .PLUS(nd_aib31_ch2_x0y0),
    .MINUS(m0_ch2_aib[31])
   );

  aliasv xaliasv30_ch2 (
    .PLUS(nd_aib30_ch2_x0y0),
    .MINUS(m0_ch2_aib[30])
   );

  aliasv xaliasv29_ch2 (
    .PLUS(nd_aib29_ch2_x0y0),
    .MINUS(m0_ch2_aib[29])
   );

  aliasv xaliasv28_ch2 (
    .PLUS(nd_aib28_ch2_x0y0),
    .MINUS(m0_ch2_aib[28])
   );

  aliasv xaliasv27_ch2 (
    .PLUS(nd_aib27_ch2_x0y0),
    .MINUS(m0_ch2_aib[27])
   );

  aliasv xaliasv26_ch2 (
    .PLUS(nd_aib26_ch2_x0y0),
    .MINUS(m0_ch2_aib[26])
   );

  aliasv xaliasv25_ch2 (
    .PLUS(nd_aib25_ch2_x0y0),
    .MINUS(m0_ch2_aib[25])
   );

  aliasv xaliasv24_ch2 (
    .PLUS(nd_aib24_ch2_x0y0),
    .MINUS(m0_ch2_aib[24])
   );

  aliasv xaliasv23_ch2 (
    .PLUS(nd_aib23_ch2_x0y0),
    .MINUS(m0_ch2_aib[23])
   );

  aliasv xaliasv22_ch2 (
    .PLUS(nd_aib22_ch2_x0y0),
    .MINUS(m0_ch2_aib[22])
   );

  aliasv xaliasv21_ch2 (
    .PLUS(nd_aib21_ch2_x0y0),
    .MINUS(m0_ch2_aib[21])
   );

  aliasv xaliasv20_ch2 (
    .PLUS(nd_aib20_ch2_x0y0),
    .MINUS(m0_ch2_aib[20])
   );

  aliasv xaliasv19_ch2 (
    .PLUS(nd_aib19_ch2_x0y0),
    .MINUS(m0_ch2_aib[19])
   );

  aliasv xaliasv18_ch2 (
    .PLUS(nd_aib18_ch2_x0y0),
    .MINUS(m0_ch2_aib[18])
   );

  aliasv xaliasv17_ch2 (
    .PLUS(nd_aib17_ch2_x0y0),
    .MINUS(m0_ch2_aib[17])
   );

  aliasv xaliasv16_ch2 (
    .PLUS(nd_aib16_ch2_x0y0),
    .MINUS(m0_ch2_aib[16])
   );

  aliasv xaliasv15_ch2 (
    .PLUS(nd_aib15_ch2_x0y0),
    .MINUS(m0_ch2_aib[15])
   );

  aliasv xaliasv14_ch2 (
    .PLUS(nd_aib14_ch2_x0y0),
    .MINUS(m0_ch2_aib[14])
   );

  aliasv xaliasv13_ch2 (
    .PLUS(nd_aib13_ch2_x0y0),
    .MINUS(m0_ch2_aib[13])
   );

  aliasv xaliasv12_ch2 (
    .PLUS(nd_aib12_ch2_x0y0),
    .MINUS(m0_ch2_aib[12])
   );

  aliasv xaliasv11_ch2 (
    .PLUS(nd_aib11_ch2_x0y0),
    .MINUS(m0_ch2_aib[11])
   );

  aliasv xaliasv10_ch2 (
    .PLUS(nd_aib10_ch2_x0y0),
    .MINUS(m0_ch2_aib[10])
   );

  aliasv xaliasv9_ch2 (
    .PLUS(nd_aib9_ch2_x0y0),
    .MINUS(m0_ch2_aib[9])
   );

  aliasv xaliasv8_ch2 (
    .PLUS(nd_aib8_ch2_x0y0),
    .MINUS(m0_ch2_aib[8])
   );

  aliasv xaliasv7_ch2 (
    .PLUS(nd_aib7_ch2_x0y0),
    .MINUS(m0_ch2_aib[7])
   );

  aliasv xaliasv6_ch2 (
    .PLUS(nd_aib6_ch2_x0y0),
    .MINUS(m0_ch2_aib[6])
   );

  aliasv xaliasv5_ch2 (
    .PLUS(nd_aib5_ch2_x0y0),
    .MINUS(m0_ch2_aib[5])
   );

  aliasv xaliasv4_ch2 (
    .PLUS(nd_aib4_ch2_x0y0),
    .MINUS(m0_ch2_aib[4])
   );

  aliasv xaliasv3_ch2 (
    .PLUS(nd_aib3_ch2_x0y0),
    .MINUS(m0_ch2_aib[3])
   );

  aliasv xaliasv2_ch2 (
    .PLUS(nd_aib2_ch2_x0y0),
    .MINUS(m0_ch2_aib[2])
   );

  aliasv xaliasv1_ch2 (
    .PLUS(nd_aib1_ch2_x0y0),
    .MINUS(m0_ch2_aib[1])
   );

  aliasv xaliasv0_ch2 (
    .PLUS(nd_aib0_ch2_x0y0),
    .MINUS(m0_ch2_aib[0])
   );

// ## START OF  ch3 ( ##
  aliasv xaliasv95_ch3 (
    .PLUS(nd_aib95_ch3_x0y0),
    .MINUS(m0_ch3_aib[95])
   );

  aliasv xaliasv94_ch3 (
    .PLUS(nd_aib94_ch3_x0y0),
    .MINUS(m0_ch3_aib[94])
   );

  aliasv xaliasv93_ch3 (
    .PLUS(nd_aib93_ch3_x0y0),
    .MINUS(m0_ch3_aib[93])
   );

  aliasv xaliasv92_ch3 (
    .PLUS(nd_aib92_ch3_x0y0),
    .MINUS(m0_ch3_aib[92])
   );

  aliasv xaliasv91_ch3 (
    .PLUS(nd_aib91_ch3_x0y0),
    .MINUS(m0_ch3_aib[91])
   );

  aliasv xaliasv90_ch3 (
    .PLUS(nd_aib90_ch3_x0y0),
    .MINUS(m0_ch3_aib[90])
   );

  aliasv xaliasv89_ch3 (
    .PLUS(nd_aib89_ch3_x0y0),
    .MINUS(m0_ch3_aib[89])
   );

  aliasv xaliasv88_ch3 (
    .PLUS(nd_aib88_ch3_x0y0),
    .MINUS(m0_ch3_aib[88])
   );

  aliasv xaliasv87_ch3 (
    .PLUS(nd_aib87_ch3_x0y0),
    .MINUS(m0_ch3_aib[87])
   );

  aliasv xaliasv86_ch3 (
    .PLUS(nd_aib86_ch3_x0y0),
    .MINUS(m0_ch3_aib[86])
   );

  aliasv xaliasv85_ch3 (
    .PLUS(nd_aib85_ch3_x0y0),
    .MINUS(m0_ch3_aib[85])
   );

  aliasv xaliasv84_ch3 (
    .PLUS(nd_aib84_ch3_x0y0),
    .MINUS(m0_ch3_aib[84])
   );

  aliasv xaliasv83_ch3 (
    .PLUS(nd_aib83_ch3_x0y0),
    .MINUS(m0_ch3_aib[83])
   );

  aliasv xaliasv82_ch3 (
    .PLUS(nd_aib82_ch3_x0y0),
    .MINUS(m0_ch3_aib[82])
   );

  aliasv xaliasv81_ch3 (
    .PLUS(nd_aib81_ch3_x0y0),
    .MINUS(m0_ch3_aib[81])
   );

  aliasv xaliasv80_ch3 (
    .PLUS(nd_aib80_ch3_x0y0),
    .MINUS(m0_ch3_aib[80])
   );

  aliasv xaliasv79_ch3 (
    .PLUS(nd_aib79_ch3_x0y0),
    .MINUS(m0_ch3_aib[79])
   );

  aliasv xaliasv78_ch3 (
    .PLUS(nd_aib78_ch3_x0y0),
    .MINUS(m0_ch3_aib[78])
   );

  aliasv xaliasv77_ch3 (
    .PLUS(nd_aib77_ch3_x0y0),
    .MINUS(m0_ch3_aib[77])
   );

  aliasv xaliasv76_ch3 (
    .PLUS(nd_aib76_ch3_x0y0),
    .MINUS(m0_ch3_aib[76])
   );

  aliasv xaliasv75_ch3 (
    .PLUS(nd_aib75_ch3_x0y0),
    .MINUS(m0_ch3_aib[75])
   );

  aliasv xaliasv74_ch3 (
    .PLUS(nd_aib74_ch3_x0y0),
    .MINUS(m0_ch3_aib[74])
   );

  aliasv xaliasv73_ch3 (
    .PLUS(nd_aib73_ch3_x0y0),
    .MINUS(m0_ch3_aib[73])
   );

  aliasv xaliasv72_ch3 (
    .PLUS(nd_aib72_ch3_x0y0),
    .MINUS(m0_ch3_aib[72])
   );

  aliasv xaliasv71_ch3 (
    .PLUS(nd_aib71_ch3_x0y0),
    .MINUS(m0_ch3_aib[71])
   );

  aliasv xaliasv70_ch3 (
    .PLUS(nd_aib70_ch3_x0y0),
    .MINUS(m0_ch3_aib[70])
   );

  aliasv xaliasv69_ch3 (
    .PLUS(nd_aib69_ch3_x0y0),
    .MINUS(m0_ch3_aib[69])
   );

  aliasv xaliasv68_ch3 (
    .PLUS(nd_aib68_ch3_x0y0),
    .MINUS(m0_ch3_aib[68])
   );

  aliasv xaliasv67_ch3 (
    .PLUS(nd_aib67_ch3_x0y0),
    .MINUS(m0_ch3_aib[67])
   );

  aliasv xaliasv66_ch3 (
    .PLUS(nd_aib66_ch3_x0y0),
    .MINUS(m0_ch3_aib[66])
   );

  aliasv xaliasv65_ch3 (
    .PLUS(nd_aib65_ch3_x0y0),
    .MINUS(m0_ch3_aib[65])
   );

  aliasv xaliasv64_ch3 (
    .PLUS(nd_aib64_ch3_x0y0),
    .MINUS(m0_ch3_aib[64])
   );

  aliasv xaliasv63_ch3 (
    .PLUS(nd_aib63_ch3_x0y0),
    .MINUS(m0_ch3_aib[63])
   );

  aliasv xaliasv62_ch3 (
    .PLUS(nd_aib62_ch3_x0y0),
    .MINUS(m0_ch3_aib[62])
   );

  aliasv xaliasv61_ch3 (
    .PLUS(nd_aib61_ch3_x0y0),
    .MINUS(m0_ch3_aib[61])
   );

  aliasv xaliasv60_ch3 (
    .PLUS(nd_aib60_ch3_x0y0),
    .MINUS(m0_ch3_aib[60])
   );

  aliasv xaliasv59_ch3 (
    .PLUS(nd_aib59_ch3_x0y0),
    .MINUS(m0_ch3_aib[59])
   );

  aliasv xaliasv58_ch3 (
    .PLUS(nd_aib58_ch3_x0y0),
    .MINUS(m0_ch3_aib[58])
   );

  aliasv xaliasv57_ch3 (
    .PLUS(nd_aib57_ch3_x0y0),
    .MINUS(m0_ch3_aib[57])
   );

  aliasv xaliasv56_ch3 (
    .PLUS(nd_aib56_ch3_x0y0),
    .MINUS(m0_ch3_aib[56])
   );

  aliasv xaliasv55_ch3 (
    .PLUS(nd_aib55_ch3_x0y0),
    .MINUS(m0_ch3_aib[55])
   );

  aliasv xaliasv54_ch3 (
    .PLUS(nd_aib54_ch3_x0y0),
    .MINUS(m0_ch3_aib[54])
   );

  aliasv xaliasv53_ch3 (
    .PLUS(nd_aib53_ch3_x0y0),
    .MINUS(m0_ch3_aib[53])
   );

  aliasv xaliasv52_ch3 (
    .PLUS(nd_aib52_ch3_x0y0),
    .MINUS(m0_ch3_aib[52])
   );

  aliasv xaliasv51_ch3 (
    .PLUS(nd_aib51_ch3_x0y0),
    .MINUS(m0_ch3_aib[51])
   );

  aliasv xaliasv50_ch3 (
    .PLUS(nd_aib50_ch3_x0y0),
    .MINUS(m0_ch3_aib[50])
   );

  aliasv xaliasv49_ch3 (
    .PLUS(nd_aib49_ch3_x0y0),
    .MINUS(m0_ch3_aib[49])
   );

  aliasv xaliasv48_ch3 (
    .PLUS(nd_aib48_ch3_x0y0),
    .MINUS(m0_ch3_aib[48])
   );

  aliasv xaliasv47_ch3 (
    .PLUS(nd_aib47_ch3_x0y0),
    .MINUS(m0_ch3_aib[47])
   );

  aliasv xaliasv46_ch3 (
    .PLUS(nd_aib46_ch3_x0y0),
    .MINUS(m0_ch3_aib[46])
   );

  aliasv xaliasv45_ch3 (
    .PLUS(nd_aib45_ch3_x0y0),
    .MINUS(m0_ch3_aib[45])
   );

  aliasv xaliasv44_ch3 (
    .PLUS(nd_aib44_ch3_x0y0),
    .MINUS(m0_ch3_aib[44])
   );

  aliasv xaliasv43_ch3 (
    .PLUS(nd_aib43_ch3_x0y0),
    .MINUS(m0_ch3_aib[43])
   );

  aliasv xaliasv42_ch3 (
    .PLUS(nd_aib42_ch3_x0y0),
    .MINUS(m0_ch3_aib[42])
   );

  aliasv xaliasv41_ch3 (
    .PLUS(nd_aib41_ch3_x0y0),
    .MINUS(m0_ch3_aib[41])
   );

  aliasv xaliasv40_ch3 (
    .PLUS(nd_aib40_ch3_x0y0),
    .MINUS(m0_ch3_aib[40])
   );

  aliasv xaliasv39_ch3 (
    .PLUS(nd_aib39_ch3_x0y0),
    .MINUS(m0_ch3_aib[39])
   );

  aliasv xaliasv38_ch3 (
    .PLUS(nd_aib38_ch3_x0y0),
    .MINUS(m0_ch3_aib[38])
   );

  aliasv xaliasv37_ch3 (
    .PLUS(nd_aib37_ch3_x0y0),
    .MINUS(m0_ch3_aib[37])
   );

  aliasv xaliasv36_ch3 (
    .PLUS(nd_aib36_ch3_x0y0),
    .MINUS(m0_ch3_aib[36])
   );

  aliasv xaliasv35_ch3 (
    .PLUS(nd_aib35_ch3_x0y0),
    .MINUS(m0_ch3_aib[35])
   );

  aliasv xaliasv34_ch3 (
    .PLUS(nd_aib34_ch3_x0y0),
    .MINUS(m0_ch3_aib[34])
   );

  aliasv xaliasv33_ch3 (
    .PLUS(nd_aib33_ch3_x0y0),
    .MINUS(m0_ch3_aib[33])
   );

  aliasv xaliasv32_ch3 (
    .PLUS(nd_aib32_ch3_x0y0),
    .MINUS(m0_ch3_aib[32])
   );

  aliasv xaliasv31_ch3 (
    .PLUS(nd_aib31_ch3_x0y0),
    .MINUS(m0_ch3_aib[31])
   );

  aliasv xaliasv30_ch3 (
    .PLUS(nd_aib30_ch3_x0y0),
    .MINUS(m0_ch3_aib[30])
   );

  aliasv xaliasv29_ch3 (
    .PLUS(nd_aib29_ch3_x0y0),
    .MINUS(m0_ch3_aib[29])
   );

  aliasv xaliasv28_ch3 (
    .PLUS(nd_aib28_ch3_x0y0),
    .MINUS(m0_ch3_aib[28])
   );

  aliasv xaliasv27_ch3 (
    .PLUS(nd_aib27_ch3_x0y0),
    .MINUS(m0_ch3_aib[27])
   );

  aliasv xaliasv26_ch3 (
    .PLUS(nd_aib26_ch3_x0y0),
    .MINUS(m0_ch3_aib[26])
   );

  aliasv xaliasv25_ch3 (
    .PLUS(nd_aib25_ch3_x0y0),
    .MINUS(m0_ch3_aib[25])
   );

  aliasv xaliasv24_ch3 (
    .PLUS(nd_aib24_ch3_x0y0),
    .MINUS(m0_ch3_aib[24])
   );

  aliasv xaliasv23_ch3 (
    .PLUS(nd_aib23_ch3_x0y0),
    .MINUS(m0_ch3_aib[23])
   );

  aliasv xaliasv22_ch3 (
    .PLUS(nd_aib22_ch3_x0y0),
    .MINUS(m0_ch3_aib[22])
   );

  aliasv xaliasv21_ch3 (
    .PLUS(nd_aib21_ch3_x0y0),
    .MINUS(m0_ch3_aib[21])
   );

  aliasv xaliasv20_ch3 (
    .PLUS(nd_aib20_ch3_x0y0),
    .MINUS(m0_ch3_aib[20])
   );

  aliasv xaliasv19_ch3 (
    .PLUS(nd_aib19_ch3_x0y0),
    .MINUS(m0_ch3_aib[19])
   );

  aliasv xaliasv18_ch3 (
    .PLUS(nd_aib18_ch3_x0y0),
    .MINUS(m0_ch3_aib[18])
   );

  aliasv xaliasv17_ch3 (
    .PLUS(nd_aib17_ch3_x0y0),
    .MINUS(m0_ch3_aib[17])
   );

  aliasv xaliasv16_ch3 (
    .PLUS(nd_aib16_ch3_x0y0),
    .MINUS(m0_ch3_aib[16])
   );

  aliasv xaliasv15_ch3 (
    .PLUS(nd_aib15_ch3_x0y0),
    .MINUS(m0_ch3_aib[15])
   );

  aliasv xaliasv14_ch3 (
    .PLUS(nd_aib14_ch3_x0y0),
    .MINUS(m0_ch3_aib[14])
   );

  aliasv xaliasv13_ch3 (
    .PLUS(nd_aib13_ch3_x0y0),
    .MINUS(m0_ch3_aib[13])
   );

  aliasv xaliasv12_ch3 (
    .PLUS(nd_aib12_ch3_x0y0),
    .MINUS(m0_ch3_aib[12])
   );

  aliasv xaliasv11_ch3 (
    .PLUS(nd_aib11_ch3_x0y0),
    .MINUS(m0_ch3_aib[11])
   );

  aliasv xaliasv10_ch3 (
    .PLUS(nd_aib10_ch3_x0y0),
    .MINUS(m0_ch3_aib[10])
   );

  aliasv xaliasv9_ch3 (
    .PLUS(nd_aib9_ch3_x0y0),
    .MINUS(m0_ch3_aib[9])
   );

  aliasv xaliasv8_ch3 (
    .PLUS(nd_aib8_ch3_x0y0),
    .MINUS(m0_ch3_aib[8])
   );

  aliasv xaliasv7_ch3 (
    .PLUS(nd_aib7_ch3_x0y0),
    .MINUS(m0_ch3_aib[7])
   );

  aliasv xaliasv6_ch3 (
    .PLUS(nd_aib6_ch3_x0y0),
    .MINUS(m0_ch3_aib[6])
   );

  aliasv xaliasv5_ch3 (
    .PLUS(nd_aib5_ch3_x0y0),
    .MINUS(m0_ch3_aib[5])
   );

  aliasv xaliasv4_ch3 (
    .PLUS(nd_aib4_ch3_x0y0),
    .MINUS(m0_ch3_aib[4])
   );

  aliasv xaliasv3_ch3 (
    .PLUS(nd_aib3_ch3_x0y0),
    .MINUS(m0_ch3_aib[3])
   );

  aliasv xaliasv2_ch3 (
    .PLUS(nd_aib2_ch3_x0y0),
    .MINUS(m0_ch3_aib[2])
   );

  aliasv xaliasv1_ch3 (
    .PLUS(nd_aib1_ch3_x0y0),
    .MINUS(m0_ch3_aib[1])
   );

  aliasv xaliasv0_ch3 (
    .PLUS(nd_aib0_ch3_x0y0),
    .MINUS(m0_ch3_aib[0])
   );

// ## START OF  ch4 ( ##
  aliasv xaliasv95_ch4 (
    .PLUS(nd_aib95_ch4_x0y0),
    .MINUS(m0_ch4_aib[95])
   );

  aliasv xaliasv94_ch4 (
    .PLUS(nd_aib94_ch4_x0y0),
    .MINUS(m0_ch4_aib[94])
   );

  aliasv xaliasv93_ch4 (
    .PLUS(nd_aib93_ch4_x0y0),
    .MINUS(m0_ch4_aib[93])
   );

  aliasv xaliasv92_ch4 (
    .PLUS(nd_aib92_ch4_x0y0),
    .MINUS(m0_ch4_aib[92])
   );

  aliasv xaliasv91_ch4 (
    .PLUS(nd_aib91_ch4_x0y0),
    .MINUS(m0_ch4_aib[91])
   );

  aliasv xaliasv90_ch4 (
    .PLUS(nd_aib90_ch4_x0y0),
    .MINUS(m0_ch4_aib[90])
   );

  aliasv xaliasv89_ch4 (
    .PLUS(nd_aib89_ch4_x0y0),
    .MINUS(m0_ch4_aib[89])
   );

  aliasv xaliasv88_ch4 (
    .PLUS(nd_aib88_ch4_x0y0),
    .MINUS(m0_ch4_aib[88])
   );

  aliasv xaliasv87_ch4 (
    .PLUS(nd_aib87_ch4_x0y0),
    .MINUS(m0_ch4_aib[87])
   );

  aliasv xaliasv86_ch4 (
    .PLUS(nd_aib86_ch4_x0y0),
    .MINUS(m0_ch4_aib[86])
   );

  aliasv xaliasv85_ch4 (
    .PLUS(nd_aib85_ch4_x0y0),
    .MINUS(m0_ch4_aib[85])
   );

  aliasv xaliasv84_ch4 (
    .PLUS(nd_aib84_ch4_x0y0),
    .MINUS(m0_ch4_aib[84])
   );

  aliasv xaliasv83_ch4 (
    .PLUS(nd_aib83_ch4_x0y0),
    .MINUS(m0_ch4_aib[83])
   );

  aliasv xaliasv82_ch4 (
    .PLUS(nd_aib82_ch4_x0y0),
    .MINUS(m0_ch4_aib[82])
   );

  aliasv xaliasv81_ch4 (
    .PLUS(nd_aib81_ch4_x0y0),
    .MINUS(m0_ch4_aib[81])
   );

  aliasv xaliasv80_ch4 (
    .PLUS(nd_aib80_ch4_x0y0),
    .MINUS(m0_ch4_aib[80])
   );

  aliasv xaliasv79_ch4 (
    .PLUS(nd_aib79_ch4_x0y0),
    .MINUS(m0_ch4_aib[79])
   );

  aliasv xaliasv78_ch4 (
    .PLUS(nd_aib78_ch4_x0y0),
    .MINUS(m0_ch4_aib[78])
   );

  aliasv xaliasv77_ch4 (
    .PLUS(nd_aib77_ch4_x0y0),
    .MINUS(m0_ch4_aib[77])
   );

  aliasv xaliasv76_ch4 (
    .PLUS(nd_aib76_ch4_x0y0),
    .MINUS(m0_ch4_aib[76])
   );

  aliasv xaliasv75_ch4 (
    .PLUS(nd_aib75_ch4_x0y0),
    .MINUS(m0_ch4_aib[75])
   );

  aliasv xaliasv74_ch4 (
    .PLUS(nd_aib74_ch4_x0y0),
    .MINUS(m0_ch4_aib[74])
   );

  aliasv xaliasv73_ch4 (
    .PLUS(nd_aib73_ch4_x0y0),
    .MINUS(m0_ch4_aib[73])
   );

  aliasv xaliasv72_ch4 (
    .PLUS(nd_aib72_ch4_x0y0),
    .MINUS(m0_ch4_aib[72])
   );

  aliasv xaliasv71_ch4 (
    .PLUS(nd_aib71_ch4_x0y0),
    .MINUS(m0_ch4_aib[71])
   );

  aliasv xaliasv70_ch4 (
    .PLUS(nd_aib70_ch4_x0y0),
    .MINUS(m0_ch4_aib[70])
   );

  aliasv xaliasv69_ch4 (
    .PLUS(nd_aib69_ch4_x0y0),
    .MINUS(m0_ch4_aib[69])
   );

  aliasv xaliasv68_ch4 (
    .PLUS(nd_aib68_ch4_x0y0),
    .MINUS(m0_ch4_aib[68])
   );

  aliasv xaliasv67_ch4 (
    .PLUS(nd_aib67_ch4_x0y0),
    .MINUS(m0_ch4_aib[67])
   );

  aliasv xaliasv66_ch4 (
    .PLUS(nd_aib66_ch4_x0y0),
    .MINUS(m0_ch4_aib[66])
   );

  aliasv xaliasv65_ch4 (
    .PLUS(nd_aib65_ch4_x0y0),
    .MINUS(m0_ch4_aib[65])
   );

  aliasv xaliasv64_ch4 (
    .PLUS(nd_aib64_ch4_x0y0),
    .MINUS(m0_ch4_aib[64])
   );

  aliasv xaliasv63_ch4 (
    .PLUS(nd_aib63_ch4_x0y0),
    .MINUS(m0_ch4_aib[63])
   );

  aliasv xaliasv62_ch4 (
    .PLUS(nd_aib62_ch4_x0y0),
    .MINUS(m0_ch4_aib[62])
   );

  aliasv xaliasv61_ch4 (
    .PLUS(nd_aib61_ch4_x0y0),
    .MINUS(m0_ch4_aib[61])
   );

  aliasv xaliasv60_ch4 (
    .PLUS(nd_aib60_ch4_x0y0),
    .MINUS(m0_ch4_aib[60])
   );

  aliasv xaliasv59_ch4 (
    .PLUS(nd_aib59_ch4_x0y0),
    .MINUS(m0_ch4_aib[59])
   );

  aliasv xaliasv58_ch4 (
    .PLUS(nd_aib58_ch4_x0y0),
    .MINUS(m0_ch4_aib[58])
   );

  aliasv xaliasv57_ch4 (
    .PLUS(nd_aib57_ch4_x0y0),
    .MINUS(m0_ch4_aib[57])
   );

  aliasv xaliasv56_ch4 (
    .PLUS(nd_aib56_ch4_x0y0),
    .MINUS(m0_ch4_aib[56])
   );

  aliasv xaliasv55_ch4 (
    .PLUS(nd_aib55_ch4_x0y0),
    .MINUS(m0_ch4_aib[55])
   );

  aliasv xaliasv54_ch4 (
    .PLUS(nd_aib54_ch4_x0y0),
    .MINUS(m0_ch4_aib[54])
   );

  aliasv xaliasv53_ch4 (
    .PLUS(nd_aib53_ch4_x0y0),
    .MINUS(m0_ch4_aib[53])
   );

  aliasv xaliasv52_ch4 (
    .PLUS(nd_aib52_ch4_x0y0),
    .MINUS(m0_ch4_aib[52])
   );

  aliasv xaliasv51_ch4 (
    .PLUS(nd_aib51_ch4_x0y0),
    .MINUS(m0_ch4_aib[51])
   );

  aliasv xaliasv50_ch4 (
    .PLUS(nd_aib50_ch4_x0y0),
    .MINUS(m0_ch4_aib[50])
   );

  aliasv xaliasv49_ch4 (
    .PLUS(nd_aib49_ch4_x0y0),
    .MINUS(m0_ch4_aib[49])
   );

  aliasv xaliasv48_ch4 (
    .PLUS(nd_aib48_ch4_x0y0),
    .MINUS(m0_ch4_aib[48])
   );

  aliasv xaliasv47_ch4 (
    .PLUS(nd_aib47_ch4_x0y0),
    .MINUS(m0_ch4_aib[47])
   );

  aliasv xaliasv46_ch4 (
    .PLUS(nd_aib46_ch4_x0y0),
    .MINUS(m0_ch4_aib[46])
   );

  aliasv xaliasv45_ch4 (
    .PLUS(nd_aib45_ch4_x0y0),
    .MINUS(m0_ch4_aib[45])
   );

  aliasv xaliasv44_ch4 (
    .PLUS(nd_aib44_ch4_x0y0),
    .MINUS(m0_ch4_aib[44])
   );

  aliasv xaliasv43_ch4 (
    .PLUS(nd_aib43_ch4_x0y0),
    .MINUS(m0_ch4_aib[43])
   );

  aliasv xaliasv42_ch4 (
    .PLUS(nd_aib42_ch4_x0y0),
    .MINUS(m0_ch4_aib[42])
   );

  aliasv xaliasv41_ch4 (
    .PLUS(nd_aib41_ch4_x0y0),
    .MINUS(m0_ch4_aib[41])
   );

  aliasv xaliasv40_ch4 (
    .PLUS(nd_aib40_ch4_x0y0),
    .MINUS(m0_ch4_aib[40])
   );

  aliasv xaliasv39_ch4 (
    .PLUS(nd_aib39_ch4_x0y0),
    .MINUS(m0_ch4_aib[39])
   );

  aliasv xaliasv38_ch4 (
    .PLUS(nd_aib38_ch4_x0y0),
    .MINUS(m0_ch4_aib[38])
   );

  aliasv xaliasv37_ch4 (
    .PLUS(nd_aib37_ch4_x0y0),
    .MINUS(m0_ch4_aib[37])
   );

  aliasv xaliasv36_ch4 (
    .PLUS(nd_aib36_ch4_x0y0),
    .MINUS(m0_ch4_aib[36])
   );

  aliasv xaliasv35_ch4 (
    .PLUS(nd_aib35_ch4_x0y0),
    .MINUS(m0_ch4_aib[35])
   );

  aliasv xaliasv34_ch4 (
    .PLUS(nd_aib34_ch4_x0y0),
    .MINUS(m0_ch4_aib[34])
   );

  aliasv xaliasv33_ch4 (
    .PLUS(nd_aib33_ch4_x0y0),
    .MINUS(m0_ch4_aib[33])
   );

  aliasv xaliasv32_ch4 (
    .PLUS(nd_aib32_ch4_x0y0),
    .MINUS(m0_ch4_aib[32])
   );

  aliasv xaliasv31_ch4 (
    .PLUS(nd_aib31_ch4_x0y0),
    .MINUS(m0_ch4_aib[31])
   );

  aliasv xaliasv30_ch4 (
    .PLUS(nd_aib30_ch4_x0y0),
    .MINUS(m0_ch4_aib[30])
   );

  aliasv xaliasv29_ch4 (
    .PLUS(nd_aib29_ch4_x0y0),
    .MINUS(m0_ch4_aib[29])
   );

  aliasv xaliasv28_ch4 (
    .PLUS(nd_aib28_ch4_x0y0),
    .MINUS(m0_ch4_aib[28])
   );

  aliasv xaliasv27_ch4 (
    .PLUS(nd_aib27_ch4_x0y0),
    .MINUS(m0_ch4_aib[27])
   );

  aliasv xaliasv26_ch4 (
    .PLUS(nd_aib26_ch4_x0y0),
    .MINUS(m0_ch4_aib[26])
   );

  aliasv xaliasv25_ch4 (
    .PLUS(nd_aib25_ch4_x0y0),
    .MINUS(m0_ch4_aib[25])
   );

  aliasv xaliasv24_ch4 (
    .PLUS(nd_aib24_ch4_x0y0),
    .MINUS(m0_ch4_aib[24])
   );

  aliasv xaliasv23_ch4 (
    .PLUS(nd_aib23_ch4_x0y0),
    .MINUS(m0_ch4_aib[23])
   );

  aliasv xaliasv22_ch4 (
    .PLUS(nd_aib22_ch4_x0y0),
    .MINUS(m0_ch4_aib[22])
   );

  aliasv xaliasv21_ch4 (
    .PLUS(nd_aib21_ch4_x0y0),
    .MINUS(m0_ch4_aib[21])
   );

  aliasv xaliasv20_ch4 (
    .PLUS(nd_aib20_ch4_x0y0),
    .MINUS(m0_ch4_aib[20])
   );

  aliasv xaliasv19_ch4 (
    .PLUS(nd_aib19_ch4_x0y0),
    .MINUS(m0_ch4_aib[19])
   );

  aliasv xaliasv18_ch4 (
    .PLUS(nd_aib18_ch4_x0y0),
    .MINUS(m0_ch4_aib[18])
   );

  aliasv xaliasv17_ch4 (
    .PLUS(nd_aib17_ch4_x0y0),
    .MINUS(m0_ch4_aib[17])
   );

  aliasv xaliasv16_ch4 (
    .PLUS(nd_aib16_ch4_x0y0),
    .MINUS(m0_ch4_aib[16])
   );

  aliasv xaliasv15_ch4 (
    .PLUS(nd_aib15_ch4_x0y0),
    .MINUS(m0_ch4_aib[15])
   );

  aliasv xaliasv14_ch4 (
    .PLUS(nd_aib14_ch4_x0y0),
    .MINUS(m0_ch4_aib[14])
   );

  aliasv xaliasv13_ch4 (
    .PLUS(nd_aib13_ch4_x0y0),
    .MINUS(m0_ch4_aib[13])
   );

  aliasv xaliasv12_ch4 (
    .PLUS(nd_aib12_ch4_x0y0),
    .MINUS(m0_ch4_aib[12])
   );

  aliasv xaliasv11_ch4 (
    .PLUS(nd_aib11_ch4_x0y0),
    .MINUS(m0_ch4_aib[11])
   );

  aliasv xaliasv10_ch4 (
    .PLUS(nd_aib10_ch4_x0y0),
    .MINUS(m0_ch4_aib[10])
   );

  aliasv xaliasv9_ch4 (
    .PLUS(nd_aib9_ch4_x0y0),
    .MINUS(m0_ch4_aib[9])
   );

  aliasv xaliasv8_ch4 (
    .PLUS(nd_aib8_ch4_x0y0),
    .MINUS(m0_ch4_aib[8])
   );

  aliasv xaliasv7_ch4 (
    .PLUS(nd_aib7_ch4_x0y0),
    .MINUS(m0_ch4_aib[7])
   );

  aliasv xaliasv6_ch4 (
    .PLUS(nd_aib6_ch4_x0y0),
    .MINUS(m0_ch4_aib[6])
   );

  aliasv xaliasv5_ch4 (
    .PLUS(nd_aib5_ch4_x0y0),
    .MINUS(m0_ch4_aib[5])
   );

  aliasv xaliasv4_ch4 (
    .PLUS(nd_aib4_ch4_x0y0),
    .MINUS(m0_ch4_aib[4])
   );

  aliasv xaliasv3_ch4 (
    .PLUS(nd_aib3_ch4_x0y0),
    .MINUS(m0_ch4_aib[3])
   );

  aliasv xaliasv2_ch4 (
    .PLUS(nd_aib2_ch4_x0y0),
    .MINUS(m0_ch4_aib[2])
   );

  aliasv xaliasv1_ch4 (
    .PLUS(nd_aib1_ch4_x0y0),
    .MINUS(m0_ch4_aib[1])
   );

  aliasv xaliasv0_ch4 (
    .PLUS(nd_aib0_ch4_x0y0),
    .MINUS(m0_ch4_aib[0])
   );

// ## START OF  ch5 ( ##
  aliasv xaliasv95_ch5 (
    .PLUS(nd_aib95_ch5_x0y0),
    .MINUS(m0_ch5_aib[95])
   );

  aliasv xaliasv94_ch5 (
    .PLUS(nd_aib94_ch5_x0y0),
    .MINUS(m0_ch5_aib[94])
   );

  aliasv xaliasv93_ch5 (
    .PLUS(nd_aib93_ch5_x0y0),
    .MINUS(m0_ch5_aib[93])
   );

  aliasv xaliasv92_ch5 (
    .PLUS(nd_aib92_ch5_x0y0),
    .MINUS(m0_ch5_aib[92])
   );

  aliasv xaliasv91_ch5 (
    .PLUS(nd_aib91_ch5_x0y0),
    .MINUS(m0_ch5_aib[91])
   );

  aliasv xaliasv90_ch5 (
    .PLUS(nd_aib90_ch5_x0y0),
    .MINUS(m0_ch5_aib[90])
   );

  aliasv xaliasv89_ch5 (
    .PLUS(nd_aib89_ch5_x0y0),
    .MINUS(m0_ch5_aib[89])
   );

  aliasv xaliasv88_ch5 (
    .PLUS(nd_aib88_ch5_x0y0),
    .MINUS(m0_ch5_aib[88])
   );

  aliasv xaliasv87_ch5 (
    .PLUS(nd_aib87_ch5_x0y0),
    .MINUS(m0_ch5_aib[87])
   );

  aliasv xaliasv86_ch5 (
    .PLUS(nd_aib86_ch5_x0y0),
    .MINUS(m0_ch5_aib[86])
   );

  aliasv xaliasv85_ch5 (
    .PLUS(nd_aib85_ch5_x0y0),
    .MINUS(m0_ch5_aib[85])
   );

  aliasv xaliasv84_ch5 (
    .PLUS(nd_aib84_ch5_x0y0),
    .MINUS(m0_ch5_aib[84])
   );

  aliasv xaliasv83_ch5 (
    .PLUS(nd_aib83_ch5_x0y0),
    .MINUS(m0_ch5_aib[83])
   );

  aliasv xaliasv82_ch5 (
    .PLUS(nd_aib82_ch5_x0y0),
    .MINUS(m0_ch5_aib[82])
   );

  aliasv xaliasv81_ch5 (
    .PLUS(nd_aib81_ch5_x0y0),
    .MINUS(m0_ch5_aib[81])
   );

  aliasv xaliasv80_ch5 (
    .PLUS(nd_aib80_ch5_x0y0),
    .MINUS(m0_ch5_aib[80])
   );

  aliasv xaliasv79_ch5 (
    .PLUS(nd_aib79_ch5_x0y0),
    .MINUS(m0_ch5_aib[79])
   );

  aliasv xaliasv78_ch5 (
    .PLUS(nd_aib78_ch5_x0y0),
    .MINUS(m0_ch5_aib[78])
   );

  aliasv xaliasv77_ch5 (
    .PLUS(nd_aib77_ch5_x0y0),
    .MINUS(m0_ch5_aib[77])
   );

  aliasv xaliasv76_ch5 (
    .PLUS(nd_aib76_ch5_x0y0),
    .MINUS(m0_ch5_aib[76])
   );

  aliasv xaliasv75_ch5 (
    .PLUS(nd_aib75_ch5_x0y0),
    .MINUS(m0_ch5_aib[75])
   );

  aliasv xaliasv74_ch5 (
    .PLUS(nd_aib74_ch5_x0y0),
    .MINUS(m0_ch5_aib[74])
   );

  aliasv xaliasv73_ch5 (
    .PLUS(nd_aib73_ch5_x0y0),
    .MINUS(m0_ch5_aib[73])
   );

  aliasv xaliasv72_ch5 (
    .PLUS(nd_aib72_ch5_x0y0),
    .MINUS(m0_ch5_aib[72])
   );

  aliasv xaliasv71_ch5 (
    .PLUS(nd_aib71_ch5_x0y0),
    .MINUS(m0_ch5_aib[71])
   );

  aliasv xaliasv70_ch5 (
    .PLUS(nd_aib70_ch5_x0y0),
    .MINUS(m0_ch5_aib[70])
   );

  aliasv xaliasv69_ch5 (
    .PLUS(nd_aib69_ch5_x0y0),
    .MINUS(m0_ch5_aib[69])
   );

  aliasv xaliasv68_ch5 (
    .PLUS(nd_aib68_ch5_x0y0),
    .MINUS(m0_ch5_aib[68])
   );

  aliasv xaliasv67_ch5 (
    .PLUS(nd_aib67_ch5_x0y0),
    .MINUS(m0_ch5_aib[67])
   );

  aliasv xaliasv66_ch5 (
    .PLUS(nd_aib66_ch5_x0y0),
    .MINUS(m0_ch5_aib[66])
   );

  aliasv xaliasv65_ch5 (
    .PLUS(nd_aib65_ch5_x0y0),
    .MINUS(m0_ch5_aib[65])
   );

  aliasv xaliasv64_ch5 (
    .PLUS(nd_aib64_ch5_x0y0),
    .MINUS(m0_ch5_aib[64])
   );

  aliasv xaliasv63_ch5 (
    .PLUS(nd_aib63_ch5_x0y0),
    .MINUS(m0_ch5_aib[63])
   );

  aliasv xaliasv62_ch5 (
    .PLUS(nd_aib62_ch5_x0y0),
    .MINUS(m0_ch5_aib[62])
   );

  aliasv xaliasv61_ch5 (
    .PLUS(nd_aib61_ch5_x0y0),
    .MINUS(m0_ch5_aib[61])
   );

  aliasv xaliasv60_ch5 (
    .PLUS(nd_aib60_ch5_x0y0),
    .MINUS(m0_ch5_aib[60])
   );

  aliasv xaliasv59_ch5 (
    .PLUS(nd_aib59_ch5_x0y0),
    .MINUS(m0_ch5_aib[59])
   );

  aliasv xaliasv58_ch5 (
    .PLUS(nd_aib58_ch5_x0y0),
    .MINUS(m0_ch5_aib[58])
   );

  aliasv xaliasv57_ch5 (
    .PLUS(nd_aib57_ch5_x0y0),
    .MINUS(m0_ch5_aib[57])
   );

  aliasv xaliasv56_ch5 (
    .PLUS(nd_aib56_ch5_x0y0),
    .MINUS(m0_ch5_aib[56])
   );

  aliasv xaliasv55_ch5 (
    .PLUS(nd_aib55_ch5_x0y0),
    .MINUS(m0_ch5_aib[55])
   );

  aliasv xaliasv54_ch5 (
    .PLUS(nd_aib54_ch5_x0y0),
    .MINUS(m0_ch5_aib[54])
   );

  aliasv xaliasv53_ch5 (
    .PLUS(nd_aib53_ch5_x0y0),
    .MINUS(m0_ch5_aib[53])
   );

  aliasv xaliasv52_ch5 (
    .PLUS(nd_aib52_ch5_x0y0),
    .MINUS(m0_ch5_aib[52])
   );

  aliasv xaliasv51_ch5 (
    .PLUS(nd_aib51_ch5_x0y0),
    .MINUS(m0_ch5_aib[51])
   );

  aliasv xaliasv50_ch5 (
    .PLUS(nd_aib50_ch5_x0y0),
    .MINUS(m0_ch5_aib[50])
   );

  aliasv xaliasv49_ch5 (
    .PLUS(nd_aib49_ch5_x0y0),
    .MINUS(m0_ch5_aib[49])
   );

  aliasv xaliasv48_ch5 (
    .PLUS(nd_aib48_ch5_x0y0),
    .MINUS(m0_ch5_aib[48])
   );

  aliasv xaliasv47_ch5 (
    .PLUS(nd_aib47_ch5_x0y0),
    .MINUS(m0_ch5_aib[47])
   );

  aliasv xaliasv46_ch5 (
    .PLUS(nd_aib46_ch5_x0y0),
    .MINUS(m0_ch5_aib[46])
   );

  aliasv xaliasv45_ch5 (
    .PLUS(nd_aib45_ch5_x0y0),
    .MINUS(m0_ch5_aib[45])
   );

  aliasv xaliasv44_ch5 (
    .PLUS(nd_aib44_ch5_x0y0),
    .MINUS(m0_ch5_aib[44])
   );

  aliasv xaliasv43_ch5 (
    .PLUS(nd_aib43_ch5_x0y0),
    .MINUS(m0_ch5_aib[43])
   );

  aliasv xaliasv42_ch5 (
    .PLUS(nd_aib42_ch5_x0y0),
    .MINUS(m0_ch5_aib[42])
   );

  aliasv xaliasv41_ch5 (
    .PLUS(nd_aib41_ch5_x0y0),
    .MINUS(m0_ch5_aib[41])
   );

  aliasv xaliasv40_ch5 (
    .PLUS(nd_aib40_ch5_x0y0),
    .MINUS(m0_ch5_aib[40])
   );

  aliasv xaliasv39_ch5 (
    .PLUS(nd_aib39_ch5_x0y0),
    .MINUS(m0_ch5_aib[39])
   );

  aliasv xaliasv38_ch5 (
    .PLUS(nd_aib38_ch5_x0y0),
    .MINUS(m0_ch5_aib[38])
   );

  aliasv xaliasv37_ch5 (
    .PLUS(nd_aib37_ch5_x0y0),
    .MINUS(m0_ch5_aib[37])
   );

  aliasv xaliasv36_ch5 (
    .PLUS(nd_aib36_ch5_x0y0),
    .MINUS(m0_ch5_aib[36])
   );

  aliasv xaliasv35_ch5 (
    .PLUS(nd_aib35_ch5_x0y0),
    .MINUS(m0_ch5_aib[35])
   );

  aliasv xaliasv34_ch5 (
    .PLUS(nd_aib34_ch5_x0y0),
    .MINUS(m0_ch5_aib[34])
   );

  aliasv xaliasv33_ch5 (
    .PLUS(nd_aib33_ch5_x0y0),
    .MINUS(m0_ch5_aib[33])
   );

  aliasv xaliasv32_ch5 (
    .PLUS(nd_aib32_ch5_x0y0),
    .MINUS(m0_ch5_aib[32])
   );

  aliasv xaliasv31_ch5 (
    .PLUS(nd_aib31_ch5_x0y0),
    .MINUS(m0_ch5_aib[31])
   );

  aliasv xaliasv30_ch5 (
    .PLUS(nd_aib30_ch5_x0y0),
    .MINUS(m0_ch5_aib[30])
   );

  aliasv xaliasv29_ch5 (
    .PLUS(nd_aib29_ch5_x0y0),
    .MINUS(m0_ch5_aib[29])
   );

  aliasv xaliasv28_ch5 (
    .PLUS(nd_aib28_ch5_x0y0),
    .MINUS(m0_ch5_aib[28])
   );

  aliasv xaliasv27_ch5 (
    .PLUS(nd_aib27_ch5_x0y0),
    .MINUS(m0_ch5_aib[27])
   );

  aliasv xaliasv26_ch5 (
    .PLUS(nd_aib26_ch5_x0y0),
    .MINUS(m0_ch5_aib[26])
   );

  aliasv xaliasv25_ch5 (
    .PLUS(nd_aib25_ch5_x0y0),
    .MINUS(m0_ch5_aib[25])
   );

  aliasv xaliasv24_ch5 (
    .PLUS(nd_aib24_ch5_x0y0),
    .MINUS(m0_ch5_aib[24])
   );

  aliasv xaliasv23_ch5 (
    .PLUS(nd_aib23_ch5_x0y0),
    .MINUS(m0_ch5_aib[23])
   );

  aliasv xaliasv22_ch5 (
    .PLUS(nd_aib22_ch5_x0y0),
    .MINUS(m0_ch5_aib[22])
   );

  aliasv xaliasv21_ch5 (
    .PLUS(nd_aib21_ch5_x0y0),
    .MINUS(m0_ch5_aib[21])
   );

  aliasv xaliasv20_ch5 (
    .PLUS(nd_aib20_ch5_x0y0),
    .MINUS(m0_ch5_aib[20])
   );

  aliasv xaliasv19_ch5 (
    .PLUS(nd_aib19_ch5_x0y0),
    .MINUS(m0_ch5_aib[19])
   );

  aliasv xaliasv18_ch5 (
    .PLUS(nd_aib18_ch5_x0y0),
    .MINUS(m0_ch5_aib[18])
   );

  aliasv xaliasv17_ch5 (
    .PLUS(nd_aib17_ch5_x0y0),
    .MINUS(m0_ch5_aib[17])
   );

  aliasv xaliasv16_ch5 (
    .PLUS(nd_aib16_ch5_x0y0),
    .MINUS(m0_ch5_aib[16])
   );

  aliasv xaliasv15_ch5 (
    .PLUS(nd_aib15_ch5_x0y0),
    .MINUS(m0_ch5_aib[15])
   );

  aliasv xaliasv14_ch5 (
    .PLUS(nd_aib14_ch5_x0y0),
    .MINUS(m0_ch5_aib[14])
   );

  aliasv xaliasv13_ch5 (
    .PLUS(nd_aib13_ch5_x0y0),
    .MINUS(m0_ch5_aib[13])
   );

  aliasv xaliasv12_ch5 (
    .PLUS(nd_aib12_ch5_x0y0),
    .MINUS(m0_ch5_aib[12])
   );

  aliasv xaliasv11_ch5 (
    .PLUS(nd_aib11_ch5_x0y0),
    .MINUS(m0_ch5_aib[11])
   );

  aliasv xaliasv10_ch5 (
    .PLUS(nd_aib10_ch5_x0y0),
    .MINUS(m0_ch5_aib[10])
   );

  aliasv xaliasv9_ch5 (
    .PLUS(nd_aib9_ch5_x0y0),
    .MINUS(m0_ch5_aib[9])
   );

  aliasv xaliasv8_ch5 (
    .PLUS(nd_aib8_ch5_x0y0),
    .MINUS(m0_ch5_aib[8])
   );

  aliasv xaliasv7_ch5 (
    .PLUS(nd_aib7_ch5_x0y0),
    .MINUS(m0_ch5_aib[7])
   );

  aliasv xaliasv6_ch5 (
    .PLUS(nd_aib6_ch5_x0y0),
    .MINUS(m0_ch5_aib[6])
   );

  aliasv xaliasv5_ch5 (
    .PLUS(nd_aib5_ch5_x0y0),
    .MINUS(m0_ch5_aib[5])
   );

  aliasv xaliasv4_ch5 (
    .PLUS(nd_aib4_ch5_x0y0),
    .MINUS(m0_ch5_aib[4])
   );

  aliasv xaliasv3_ch5 (
    .PLUS(nd_aib3_ch5_x0y0),
    .MINUS(m0_ch5_aib[3])
   );

  aliasv xaliasv2_ch5 (
    .PLUS(nd_aib2_ch5_x0y0),
    .MINUS(m0_ch5_aib[2])
   );

  aliasv xaliasv1_ch5 (
    .PLUS(nd_aib1_ch5_x0y0),
    .MINUS(m0_ch5_aib[1])
   );

  aliasv xaliasv0_ch5 (
    .PLUS(nd_aib0_ch5_x0y0),
    .MINUS(m0_ch5_aib[0])
   );

// ## START OF  ch6 ( ##
  aliasv xaliasv95_ch6 (
    .PLUS(nd_aib95_ch0_x0y1),
    .MINUS(m1_ch0_aib[95])
   );

  aliasv xaliasv94_ch6 (
    .PLUS(nd_aib94_ch0_x0y1),
    .MINUS(m1_ch0_aib[94])
   );

  aliasv xaliasv93_ch6 (
    .PLUS(nd_aib93_ch0_x0y1),
    .MINUS(m1_ch0_aib[93])
   );

  aliasv xaliasv92_ch6 (
    .PLUS(nd_aib92_ch0_x0y1),
    .MINUS(m1_ch0_aib[92])
   );

  aliasv xaliasv91_ch6 (
    .PLUS(nd_aib91_ch0_x0y1),
    .MINUS(m1_ch0_aib[91])
   );

  aliasv xaliasv90_ch6 (
    .PLUS(nd_aib90_ch0_x0y1),
    .MINUS(m1_ch0_aib[90])
   );

  aliasv xaliasv89_ch6 (
    .PLUS(nd_aib89_ch0_x0y1),
    .MINUS(m1_ch0_aib[89])
   );

  aliasv xaliasv88_ch6 (
    .PLUS(nd_aib88_ch0_x0y1),
    .MINUS(m1_ch0_aib[88])
   );

  aliasv xaliasv87_ch6 (
    .PLUS(nd_aib87_ch0_x0y1),
    .MINUS(m1_ch0_aib[87])
   );

  aliasv xaliasv86_ch6 (
    .PLUS(nd_aib86_ch0_x0y1),
    .MINUS(m1_ch0_aib[86])
   );

  aliasv xaliasv85_ch6 (
    .PLUS(nd_aib85_ch0_x0y1),
    .MINUS(m1_ch0_aib[85])
   );

  aliasv xaliasv84_ch6 (
    .PLUS(nd_aib84_ch0_x0y1),
    .MINUS(m1_ch0_aib[84])
   );

  aliasv xaliasv83_ch6 (
    .PLUS(nd_aib83_ch0_x0y1),
    .MINUS(m1_ch0_aib[83])
   );

  aliasv xaliasv82_ch6 (
    .PLUS(nd_aib82_ch0_x0y1),
    .MINUS(m1_ch0_aib[82])
   );

  aliasv xaliasv81_ch6 (
    .PLUS(nd_aib81_ch0_x0y1),
    .MINUS(m1_ch0_aib[81])
   );

  aliasv xaliasv80_ch6 (
    .PLUS(nd_aib80_ch0_x0y1),
    .MINUS(m1_ch0_aib[80])
   );

  aliasv xaliasv79_ch6 (
    .PLUS(nd_aib79_ch0_x0y1),
    .MINUS(m1_ch0_aib[79])
   );

  aliasv xaliasv78_ch6 (
    .PLUS(nd_aib78_ch0_x0y1),
    .MINUS(m1_ch0_aib[78])
   );

  aliasv xaliasv77_ch6 (
    .PLUS(nd_aib77_ch0_x0y1),
    .MINUS(m1_ch0_aib[77])
   );

  aliasv xaliasv76_ch6 (
    .PLUS(nd_aib76_ch0_x0y1),
    .MINUS(m1_ch0_aib[76])
   );

  aliasv xaliasv75_ch6 (
    .PLUS(nd_aib75_ch0_x0y1),
    .MINUS(m1_ch0_aib[75])
   );

  aliasv xaliasv74_ch6 (
    .PLUS(nd_aib74_ch0_x0y1),
    .MINUS(m1_ch0_aib[74])
   );

  aliasv xaliasv73_ch6 (
    .PLUS(nd_aib73_ch0_x0y1),
    .MINUS(m1_ch0_aib[73])
   );

  aliasv xaliasv72_ch6 (
    .PLUS(nd_aib72_ch0_x0y1),
    .MINUS(m1_ch0_aib[72])
   );

  aliasv xaliasv71_ch6 (
    .PLUS(nd_aib71_ch0_x0y1),
    .MINUS(m1_ch0_aib[71])
   );

  aliasv xaliasv70_ch6 (
    .PLUS(nd_aib70_ch0_x0y1),
    .MINUS(m1_ch0_aib[70])
   );

  aliasv xaliasv69_ch6 (
    .PLUS(nd_aib69_ch0_x0y1),
    .MINUS(m1_ch0_aib[69])
   );

  aliasv xaliasv68_ch6 (
    .PLUS(nd_aib68_ch0_x0y1),
    .MINUS(m1_ch0_aib[68])
   );

  aliasv xaliasv67_ch6 (
    .PLUS(nd_aib67_ch0_x0y1),
    .MINUS(m1_ch0_aib[67])
   );

  aliasv xaliasv66_ch6 (
    .PLUS(nd_aib66_ch0_x0y1),
    .MINUS(m1_ch0_aib[66])
   );

  aliasv xaliasv65_ch6 (
    .PLUS(nd_aib65_ch0_x0y1),
    .MINUS(m1_ch0_aib[65])
   );

  aliasv xaliasv64_ch6 (
    .PLUS(nd_aib64_ch0_x0y1),
    .MINUS(m1_ch0_aib[64])
   );

  aliasv xaliasv63_ch6 (
    .PLUS(nd_aib63_ch0_x0y1),
    .MINUS(m1_ch0_aib[63])
   );

  aliasv xaliasv62_ch6 (
    .PLUS(nd_aib62_ch0_x0y1),
    .MINUS(m1_ch0_aib[62])
   );

  aliasv xaliasv61_ch6 (
    .PLUS(nd_aib61_ch0_x0y1),
    .MINUS(m1_ch0_aib[61])
   );

  aliasv xaliasv60_ch6 (
    .PLUS(nd_aib60_ch0_x0y1),
    .MINUS(m1_ch0_aib[60])
   );

  aliasv xaliasv59_ch6 (
    .PLUS(nd_aib59_ch0_x0y1),
    .MINUS(m1_ch0_aib[59])
   );

  aliasv xaliasv58_ch6 (
    .PLUS(nd_aib58_ch0_x0y1),
    .MINUS(m1_ch0_aib[58])
   );

  aliasv xaliasv57_ch6 (
    .PLUS(nd_aib57_ch0_x0y1),
    .MINUS(m1_ch0_aib[57])
   );

  aliasv xaliasv56_ch6 (
    .PLUS(nd_aib56_ch0_x0y1),
    .MINUS(m1_ch0_aib[56])
   );

  aliasv xaliasv55_ch6 (
    .PLUS(nd_aib55_ch0_x0y1),
    .MINUS(m1_ch0_aib[55])
   );

  aliasv xaliasv54_ch6 (
    .PLUS(nd_aib54_ch0_x0y1),
    .MINUS(m1_ch0_aib[54])
   );

  aliasv xaliasv53_ch6 (
    .PLUS(nd_aib53_ch0_x0y1),
    .MINUS(m1_ch0_aib[53])
   );

  aliasv xaliasv52_ch6 (
    .PLUS(nd_aib52_ch0_x0y1),
    .MINUS(m1_ch0_aib[52])
   );

  aliasv xaliasv51_ch6 (
    .PLUS(nd_aib51_ch0_x0y1),
    .MINUS(m1_ch0_aib[51])
   );

  aliasv xaliasv50_ch6 (
    .PLUS(nd_aib50_ch0_x0y1),
    .MINUS(m1_ch0_aib[50])
   );

  aliasv xaliasv49_ch6 (
    .PLUS(nd_aib49_ch0_x0y1),
    .MINUS(m1_ch0_aib[49])
   );

  aliasv xaliasv48_ch6 (
    .PLUS(nd_aib48_ch0_x0y1),
    .MINUS(m1_ch0_aib[48])
   );

  aliasv xaliasv47_ch6 (
    .PLUS(nd_aib47_ch0_x0y1),
    .MINUS(m1_ch0_aib[47])
   );

  aliasv xaliasv46_ch6 (
    .PLUS(nd_aib46_ch0_x0y1),
    .MINUS(m1_ch0_aib[46])
   );

  aliasv xaliasv45_ch6 (
    .PLUS(nd_aib45_ch0_x0y1),
    .MINUS(m1_ch0_aib[45])
   );

  aliasv xaliasv44_ch6 (
    .PLUS(nd_aib44_ch0_x0y1),
    .MINUS(m1_ch0_aib[44])
   );

  aliasv xaliasv43_ch6 (
    .PLUS(nd_aib43_ch0_x0y1),
    .MINUS(m1_ch0_aib[43])
   );

  aliasv xaliasv42_ch6 (
    .PLUS(nd_aib42_ch0_x0y1),
    .MINUS(m1_ch0_aib[42])
   );

  aliasv xaliasv41_ch6 (
    .PLUS(nd_aib41_ch0_x0y1),
    .MINUS(m1_ch0_aib[41])
   );

  aliasv xaliasv40_ch6 (
    .PLUS(nd_aib40_ch0_x0y1),
    .MINUS(m1_ch0_aib[40])
   );

  aliasv xaliasv39_ch6 (
    .PLUS(nd_aib39_ch0_x0y1),
    .MINUS(m1_ch0_aib[39])
   );

  aliasv xaliasv38_ch6 (
    .PLUS(nd_aib38_ch0_x0y1),
    .MINUS(m1_ch0_aib[38])
   );

  aliasv xaliasv37_ch6 (
    .PLUS(nd_aib37_ch0_x0y1),
    .MINUS(m1_ch0_aib[37])
   );

  aliasv xaliasv36_ch6 (
    .PLUS(nd_aib36_ch0_x0y1),
    .MINUS(m1_ch0_aib[36])
   );

  aliasv xaliasv35_ch6 (
    .PLUS(nd_aib35_ch0_x0y1),
    .MINUS(m1_ch0_aib[35])
   );

  aliasv xaliasv34_ch6 (
    .PLUS(nd_aib34_ch0_x0y1),
    .MINUS(m1_ch0_aib[34])
   );

  aliasv xaliasv33_ch6 (
    .PLUS(nd_aib33_ch0_x0y1),
    .MINUS(m1_ch0_aib[33])
   );

  aliasv xaliasv32_ch6 (
    .PLUS(nd_aib32_ch0_x0y1),
    .MINUS(m1_ch0_aib[32])
   );

  aliasv xaliasv31_ch6 (
    .PLUS(nd_aib31_ch0_x0y1),
    .MINUS(m1_ch0_aib[31])
   );

  aliasv xaliasv30_ch6 (
    .PLUS(nd_aib30_ch0_x0y1),
    .MINUS(m1_ch0_aib[30])
   );

  aliasv xaliasv29_ch6 (
    .PLUS(nd_aib29_ch0_x0y1),
    .MINUS(m1_ch0_aib[29])
   );

  aliasv xaliasv28_ch6 (
    .PLUS(nd_aib28_ch0_x0y1),
    .MINUS(m1_ch0_aib[28])
   );

  aliasv xaliasv27_ch6 (
    .PLUS(nd_aib27_ch0_x0y1),
    .MINUS(m1_ch0_aib[27])
   );

  aliasv xaliasv26_ch6 (
    .PLUS(nd_aib26_ch0_x0y1),
    .MINUS(m1_ch0_aib[26])
   );

  aliasv xaliasv25_ch6 (
    .PLUS(nd_aib25_ch0_x0y1),
    .MINUS(m1_ch0_aib[25])
   );

  aliasv xaliasv24_ch6 (
    .PLUS(nd_aib24_ch0_x0y1),
    .MINUS(m1_ch0_aib[24])
   );

  aliasv xaliasv23_ch6 (
    .PLUS(nd_aib23_ch0_x0y1),
    .MINUS(m1_ch0_aib[23])
   );

  aliasv xaliasv22_ch6 (
    .PLUS(nd_aib22_ch0_x0y1),
    .MINUS(m1_ch0_aib[22])
   );

  aliasv xaliasv21_ch6 (
    .PLUS(nd_aib21_ch0_x0y1),
    .MINUS(m1_ch0_aib[21])
   );

  aliasv xaliasv20_ch6 (
    .PLUS(nd_aib20_ch0_x0y1),
    .MINUS(m1_ch0_aib[20])
   );

  aliasv xaliasv19_ch6 (
    .PLUS(nd_aib19_ch0_x0y1),
    .MINUS(m1_ch0_aib[19])
   );

  aliasv xaliasv18_ch6 (
    .PLUS(nd_aib18_ch0_x0y1),
    .MINUS(m1_ch0_aib[18])
   );

  aliasv xaliasv17_ch6 (
    .PLUS(nd_aib17_ch0_x0y1),
    .MINUS(m1_ch0_aib[17])
   );

  aliasv xaliasv16_ch6 (
    .PLUS(nd_aib16_ch0_x0y1),
    .MINUS(m1_ch0_aib[16])
   );

  aliasv xaliasv15_ch6 (
    .PLUS(nd_aib15_ch0_x0y1),
    .MINUS(m1_ch0_aib[15])
   );

  aliasv xaliasv14_ch6 (
    .PLUS(nd_aib14_ch0_x0y1),
    .MINUS(m1_ch0_aib[14])
   );

  aliasv xaliasv13_ch6 (
    .PLUS(nd_aib13_ch0_x0y1),
    .MINUS(m1_ch0_aib[13])
   );

  aliasv xaliasv12_ch6 (
    .PLUS(nd_aib12_ch0_x0y1),
    .MINUS(m1_ch0_aib[12])
   );

  aliasv xaliasv11_ch6 (
    .PLUS(nd_aib11_ch0_x0y1),
    .MINUS(m1_ch0_aib[11])
   );

  aliasv xaliasv10_ch6 (
    .PLUS(nd_aib10_ch0_x0y1),
    .MINUS(m1_ch0_aib[10])
   );

  aliasv xaliasv9_ch6 (
    .PLUS(nd_aib9_ch0_x0y1),
    .MINUS(m1_ch0_aib[9])
   );

  aliasv xaliasv8_ch6 (
    .PLUS(nd_aib8_ch0_x0y1),
    .MINUS(m1_ch0_aib[8])
   );

  aliasv xaliasv7_ch6 (
    .PLUS(nd_aib7_ch0_x0y1),
    .MINUS(m1_ch0_aib[7])
   );

  aliasv xaliasv6_ch6 (
    .PLUS(nd_aib6_ch0_x0y1),
    .MINUS(m1_ch0_aib[6])
   );

  aliasv xaliasv5_ch6 (
    .PLUS(nd_aib5_ch0_x0y1),
    .MINUS(m1_ch0_aib[5])
   );

  aliasv xaliasv4_ch6 (
    .PLUS(nd_aib4_ch0_x0y1),
    .MINUS(m1_ch0_aib[4])
   );

  aliasv xaliasv3_ch6 (
    .PLUS(nd_aib3_ch0_x0y1),
    .MINUS(m1_ch0_aib[3])
   );

  aliasv xaliasv2_ch6 (
    .PLUS(nd_aib2_ch0_x0y1),
    .MINUS(m1_ch0_aib[2])
   );

  aliasv xaliasv1_ch6 (
    .PLUS(nd_aib1_ch0_x0y1),
    .MINUS(m1_ch0_aib[1])
   );

  aliasv xaliasv0_ch6 (
    .PLUS(nd_aib0_ch0_x0y1),
    .MINUS(m1_ch0_aib[0])
   );

// ## START OF  ch7 ( ##
  aliasv xaliasv95_ch7 (
    .PLUS(nd_aib95_ch1_x0y1),
    .MINUS(m1_ch1_aib[95])
   );

  aliasv xaliasv94_ch7 (
    .PLUS(nd_aib94_ch1_x0y1),
    .MINUS(m1_ch1_aib[94])
   );

  aliasv xaliasv93_ch7 (
    .PLUS(nd_aib93_ch1_x0y1),
    .MINUS(m1_ch1_aib[93])
   );

  aliasv xaliasv92_ch7 (
    .PLUS(nd_aib92_ch1_x0y1),
    .MINUS(m1_ch1_aib[92])
   );

  aliasv xaliasv91_ch7 (
    .PLUS(nd_aib91_ch1_x0y1),
    .MINUS(m1_ch1_aib[91])
   );

  aliasv xaliasv90_ch7 (
    .PLUS(nd_aib90_ch1_x0y1),
    .MINUS(m1_ch1_aib[90])
   );

  aliasv xaliasv89_ch7 (
    .PLUS(nd_aib89_ch1_x0y1),
    .MINUS(m1_ch1_aib[89])
   );

  aliasv xaliasv88_ch7 (
    .PLUS(nd_aib88_ch1_x0y1),
    .MINUS(m1_ch1_aib[88])
   );

  aliasv xaliasv87_ch7 (
    .PLUS(nd_aib87_ch1_x0y1),
    .MINUS(m1_ch1_aib[87])
   );

  aliasv xaliasv86_ch7 (
    .PLUS(nd_aib86_ch1_x0y1),
    .MINUS(m1_ch1_aib[86])
   );

  aliasv xaliasv85_ch7 (
    .PLUS(nd_aib85_ch1_x0y1),
    .MINUS(m1_ch1_aib[85])
   );

  aliasv xaliasv84_ch7 (
    .PLUS(nd_aib84_ch1_x0y1),
    .MINUS(m1_ch1_aib[84])
   );

  aliasv xaliasv83_ch7 (
    .PLUS(nd_aib83_ch1_x0y1),
    .MINUS(m1_ch1_aib[83])
   );

  aliasv xaliasv82_ch7 (
    .PLUS(nd_aib82_ch1_x0y1),
    .MINUS(m1_ch1_aib[82])
   );

  aliasv xaliasv81_ch7 (
    .PLUS(nd_aib81_ch1_x0y1),
    .MINUS(m1_ch1_aib[81])
   );

  aliasv xaliasv80_ch7 (
    .PLUS(nd_aib80_ch1_x0y1),
    .MINUS(m1_ch1_aib[80])
   );

  aliasv xaliasv79_ch7 (
    .PLUS(nd_aib79_ch1_x0y1),
    .MINUS(m1_ch1_aib[79])
   );

  aliasv xaliasv78_ch7 (
    .PLUS(nd_aib78_ch1_x0y1),
    .MINUS(m1_ch1_aib[78])
   );

  aliasv xaliasv77_ch7 (
    .PLUS(nd_aib77_ch1_x0y1),
    .MINUS(m1_ch1_aib[77])
   );

  aliasv xaliasv76_ch7 (
    .PLUS(nd_aib76_ch1_x0y1),
    .MINUS(m1_ch1_aib[76])
   );

  aliasv xaliasv75_ch7 (
    .PLUS(nd_aib75_ch1_x0y1),
    .MINUS(m1_ch1_aib[75])
   );

  aliasv xaliasv74_ch7 (
    .PLUS(nd_aib74_ch1_x0y1),
    .MINUS(m1_ch1_aib[74])
   );

  aliasv xaliasv73_ch7 (
    .PLUS(nd_aib73_ch1_x0y1),
    .MINUS(m1_ch1_aib[73])
   );

  aliasv xaliasv72_ch7 (
    .PLUS(nd_aib72_ch1_x0y1),
    .MINUS(m1_ch1_aib[72])
   );

  aliasv xaliasv71_ch7 (
    .PLUS(nd_aib71_ch1_x0y1),
    .MINUS(m1_ch1_aib[71])
   );

  aliasv xaliasv70_ch7 (
    .PLUS(nd_aib70_ch1_x0y1),
    .MINUS(m1_ch1_aib[70])
   );

  aliasv xaliasv69_ch7 (
    .PLUS(nd_aib69_ch1_x0y1),
    .MINUS(m1_ch1_aib[69])
   );

  aliasv xaliasv68_ch7 (
    .PLUS(nd_aib68_ch1_x0y1),
    .MINUS(m1_ch1_aib[68])
   );

  aliasv xaliasv67_ch7 (
    .PLUS(nd_aib67_ch1_x0y1),
    .MINUS(m1_ch1_aib[67])
   );

  aliasv xaliasv66_ch7 (
    .PLUS(nd_aib66_ch1_x0y1),
    .MINUS(m1_ch1_aib[66])
   );

  aliasv xaliasv65_ch7 (
    .PLUS(nd_aib65_ch1_x0y1),
    .MINUS(m1_ch1_aib[65])
   );

  aliasv xaliasv64_ch7 (
    .PLUS(nd_aib64_ch1_x0y1),
    .MINUS(m1_ch1_aib[64])
   );

  aliasv xaliasv63_ch7 (
    .PLUS(nd_aib63_ch1_x0y1),
    .MINUS(m1_ch1_aib[63])
   );

  aliasv xaliasv62_ch7 (
    .PLUS(nd_aib62_ch1_x0y1),
    .MINUS(m1_ch1_aib[62])
   );

  aliasv xaliasv61_ch7 (
    .PLUS(nd_aib61_ch1_x0y1),
    .MINUS(m1_ch1_aib[61])
   );

  aliasv xaliasv60_ch7 (
    .PLUS(nd_aib60_ch1_x0y1),
    .MINUS(m1_ch1_aib[60])
   );

  aliasv xaliasv59_ch7 (
    .PLUS(nd_aib59_ch1_x0y1),
    .MINUS(m1_ch1_aib[59])
   );

  aliasv xaliasv58_ch7 (
    .PLUS(nd_aib58_ch1_x0y1),
    .MINUS(m1_ch1_aib[58])
   );

  aliasv xaliasv57_ch7 (
    .PLUS(nd_aib57_ch1_x0y1),
    .MINUS(m1_ch1_aib[57])
   );

  aliasv xaliasv56_ch7 (
    .PLUS(nd_aib56_ch1_x0y1),
    .MINUS(m1_ch1_aib[56])
   );

  aliasv xaliasv55_ch7 (
    .PLUS(nd_aib55_ch1_x0y1),
    .MINUS(m1_ch1_aib[55])
   );

  aliasv xaliasv54_ch7 (
    .PLUS(nd_aib54_ch1_x0y1),
    .MINUS(m1_ch1_aib[54])
   );

  aliasv xaliasv53_ch7 (
    .PLUS(nd_aib53_ch1_x0y1),
    .MINUS(m1_ch1_aib[53])
   );

  aliasv xaliasv52_ch7 (
    .PLUS(nd_aib52_ch1_x0y1),
    .MINUS(m1_ch1_aib[52])
   );

  aliasv xaliasv51_ch7 (
    .PLUS(nd_aib51_ch1_x0y1),
    .MINUS(m1_ch1_aib[51])
   );

  aliasv xaliasv50_ch7 (
    .PLUS(nd_aib50_ch1_x0y1),
    .MINUS(m1_ch1_aib[50])
   );

  aliasv xaliasv49_ch7 (
    .PLUS(nd_aib49_ch1_x0y1),
    .MINUS(m1_ch1_aib[49])
   );

  aliasv xaliasv48_ch7 (
    .PLUS(nd_aib48_ch1_x0y1),
    .MINUS(m1_ch1_aib[48])
   );

  aliasv xaliasv47_ch7 (
    .PLUS(nd_aib47_ch1_x0y1),
    .MINUS(m1_ch1_aib[47])
   );

  aliasv xaliasv46_ch7 (
    .PLUS(nd_aib46_ch1_x0y1),
    .MINUS(m1_ch1_aib[46])
   );

  aliasv xaliasv45_ch7 (
    .PLUS(nd_aib45_ch1_x0y1),
    .MINUS(m1_ch1_aib[45])
   );

  aliasv xaliasv44_ch7 (
    .PLUS(nd_aib44_ch1_x0y1),
    .MINUS(m1_ch1_aib[44])
   );

  aliasv xaliasv43_ch7 (
    .PLUS(nd_aib43_ch1_x0y1),
    .MINUS(m1_ch1_aib[43])
   );

  aliasv xaliasv42_ch7 (
    .PLUS(nd_aib42_ch1_x0y1),
    .MINUS(m1_ch1_aib[42])
   );

  aliasv xaliasv41_ch7 (
    .PLUS(nd_aib41_ch1_x0y1),
    .MINUS(m1_ch1_aib[41])
   );

  aliasv xaliasv40_ch7 (
    .PLUS(nd_aib40_ch1_x0y1),
    .MINUS(m1_ch1_aib[40])
   );

  aliasv xaliasv39_ch7 (
    .PLUS(nd_aib39_ch1_x0y1),
    .MINUS(m1_ch1_aib[39])
   );

  aliasv xaliasv38_ch7 (
    .PLUS(nd_aib38_ch1_x0y1),
    .MINUS(m1_ch1_aib[38])
   );

  aliasv xaliasv37_ch7 (
    .PLUS(nd_aib37_ch1_x0y1),
    .MINUS(m1_ch1_aib[37])
   );

  aliasv xaliasv36_ch7 (
    .PLUS(nd_aib36_ch1_x0y1),
    .MINUS(m1_ch1_aib[36])
   );

  aliasv xaliasv35_ch7 (
    .PLUS(nd_aib35_ch1_x0y1),
    .MINUS(m1_ch1_aib[35])
   );

  aliasv xaliasv34_ch7 (
    .PLUS(nd_aib34_ch1_x0y1),
    .MINUS(m1_ch1_aib[34])
   );

  aliasv xaliasv33_ch7 (
    .PLUS(nd_aib33_ch1_x0y1),
    .MINUS(m1_ch1_aib[33])
   );

  aliasv xaliasv32_ch7 (
    .PLUS(nd_aib32_ch1_x0y1),
    .MINUS(m1_ch1_aib[32])
   );

  aliasv xaliasv31_ch7 (
    .PLUS(nd_aib31_ch1_x0y1),
    .MINUS(m1_ch1_aib[31])
   );

  aliasv xaliasv30_ch7 (
    .PLUS(nd_aib30_ch1_x0y1),
    .MINUS(m1_ch1_aib[30])
   );

  aliasv xaliasv29_ch7 (
    .PLUS(nd_aib29_ch1_x0y1),
    .MINUS(m1_ch1_aib[29])
   );

  aliasv xaliasv28_ch7 (
    .PLUS(nd_aib28_ch1_x0y1),
    .MINUS(m1_ch1_aib[28])
   );

  aliasv xaliasv27_ch7 (
    .PLUS(nd_aib27_ch1_x0y1),
    .MINUS(m1_ch1_aib[27])
   );

  aliasv xaliasv26_ch7 (
    .PLUS(nd_aib26_ch1_x0y1),
    .MINUS(m1_ch1_aib[26])
   );

  aliasv xaliasv25_ch7 (
    .PLUS(nd_aib25_ch1_x0y1),
    .MINUS(m1_ch1_aib[25])
   );

  aliasv xaliasv24_ch7 (
    .PLUS(nd_aib24_ch1_x0y1),
    .MINUS(m1_ch1_aib[24])
   );

  aliasv xaliasv23_ch7 (
    .PLUS(nd_aib23_ch1_x0y1),
    .MINUS(m1_ch1_aib[23])
   );

  aliasv xaliasv22_ch7 (
    .PLUS(nd_aib22_ch1_x0y1),
    .MINUS(m1_ch1_aib[22])
   );

  aliasv xaliasv21_ch7 (
    .PLUS(nd_aib21_ch1_x0y1),
    .MINUS(m1_ch1_aib[21])
   );

  aliasv xaliasv20_ch7 (
    .PLUS(nd_aib20_ch1_x0y1),
    .MINUS(m1_ch1_aib[20])
   );

  aliasv xaliasv19_ch7 (
    .PLUS(nd_aib19_ch1_x0y1),
    .MINUS(m1_ch1_aib[19])
   );

  aliasv xaliasv18_ch7 (
    .PLUS(nd_aib18_ch1_x0y1),
    .MINUS(m1_ch1_aib[18])
   );

  aliasv xaliasv17_ch7 (
    .PLUS(nd_aib17_ch1_x0y1),
    .MINUS(m1_ch1_aib[17])
   );

  aliasv xaliasv16_ch7 (
    .PLUS(nd_aib16_ch1_x0y1),
    .MINUS(m1_ch1_aib[16])
   );

  aliasv xaliasv15_ch7 (
    .PLUS(nd_aib15_ch1_x0y1),
    .MINUS(m1_ch1_aib[15])
   );

  aliasv xaliasv14_ch7 (
    .PLUS(nd_aib14_ch1_x0y1),
    .MINUS(m1_ch1_aib[14])
   );

  aliasv xaliasv13_ch7 (
    .PLUS(nd_aib13_ch1_x0y1),
    .MINUS(m1_ch1_aib[13])
   );

  aliasv xaliasv12_ch7 (
    .PLUS(nd_aib12_ch1_x0y1),
    .MINUS(m1_ch1_aib[12])
   );

  aliasv xaliasv11_ch7 (
    .PLUS(nd_aib11_ch1_x0y1),
    .MINUS(m1_ch1_aib[11])
   );

  aliasv xaliasv10_ch7 (
    .PLUS(nd_aib10_ch1_x0y1),
    .MINUS(m1_ch1_aib[10])
   );

  aliasv xaliasv9_ch7 (
    .PLUS(nd_aib9_ch1_x0y1),
    .MINUS(m1_ch1_aib[9])
   );

  aliasv xaliasv8_ch7 (
    .PLUS(nd_aib8_ch1_x0y1),
    .MINUS(m1_ch1_aib[8])
   );

  aliasv xaliasv7_ch7 (
    .PLUS(nd_aib7_ch1_x0y1),
    .MINUS(m1_ch1_aib[7])
   );

  aliasv xaliasv6_ch7 (
    .PLUS(nd_aib6_ch1_x0y1),
    .MINUS(m1_ch1_aib[6])
   );

  aliasv xaliasv5_ch7 (
    .PLUS(nd_aib5_ch1_x0y1),
    .MINUS(m1_ch1_aib[5])
   );

  aliasv xaliasv4_ch7 (
    .PLUS(nd_aib4_ch1_x0y1),
    .MINUS(m1_ch1_aib[4])
   );

  aliasv xaliasv3_ch7 (
    .PLUS(nd_aib3_ch1_x0y1),
    .MINUS(m1_ch1_aib[3])
   );

  aliasv xaliasv2_ch7 (
    .PLUS(nd_aib2_ch1_x0y1),
    .MINUS(m1_ch1_aib[2])
   );

  aliasv xaliasv1_ch7 (
    .PLUS(nd_aib1_ch1_x0y1),
    .MINUS(m1_ch1_aib[1])
   );

  aliasv xaliasv0_ch7 (
    .PLUS(nd_aib0_ch1_x0y1),
    .MINUS(m1_ch1_aib[0])
   );

// ## START OF  ch8 ( ##
  aliasv xaliasv95_ch8 (
    .PLUS(nd_aib95_ch2_x0y1),
    .MINUS(m1_ch2_aib[95])
   );

  aliasv xaliasv94_ch8 (
    .PLUS(nd_aib94_ch2_x0y1),
    .MINUS(m1_ch2_aib[94])
   );

  aliasv xaliasv93_ch8 (
    .PLUS(nd_aib93_ch2_x0y1),
    .MINUS(m1_ch2_aib[93])
   );

  aliasv xaliasv92_ch8 (
    .PLUS(nd_aib92_ch2_x0y1),
    .MINUS(m1_ch2_aib[92])
   );

  aliasv xaliasv91_ch8 (
    .PLUS(nd_aib91_ch2_x0y1),
    .MINUS(m1_ch2_aib[91])
   );

  aliasv xaliasv90_ch8 (
    .PLUS(nd_aib90_ch2_x0y1),
    .MINUS(m1_ch2_aib[90])
   );

  aliasv xaliasv89_ch8 (
    .PLUS(nd_aib89_ch2_x0y1),
    .MINUS(m1_ch2_aib[89])
   );

  aliasv xaliasv88_ch8 (
    .PLUS(nd_aib88_ch2_x0y1),
    .MINUS(m1_ch2_aib[88])
   );

  aliasv xaliasv87_ch8 (
    .PLUS(nd_aib87_ch2_x0y1),
    .MINUS(m1_ch2_aib[87])
   );

  aliasv xaliasv86_ch8 (
    .PLUS(nd_aib86_ch2_x0y1),
    .MINUS(m1_ch2_aib[86])
   );

  aliasv xaliasv85_ch8 (
    .PLUS(nd_aib85_ch2_x0y1),
    .MINUS(m1_ch2_aib[85])
   );

  aliasv xaliasv84_ch8 (
    .PLUS(nd_aib84_ch2_x0y1),
    .MINUS(m1_ch2_aib[84])
   );

  aliasv xaliasv83_ch8 (
    .PLUS(nd_aib83_ch2_x0y1),
    .MINUS(m1_ch2_aib[83])
   );

  aliasv xaliasv82_ch8 (
    .PLUS(nd_aib82_ch2_x0y1),
    .MINUS(m1_ch2_aib[82])
   );

  aliasv xaliasv81_ch8 (
    .PLUS(nd_aib81_ch2_x0y1),
    .MINUS(m1_ch2_aib[81])
   );

  aliasv xaliasv80_ch8 (
    .PLUS(nd_aib80_ch2_x0y1),
    .MINUS(m1_ch2_aib[80])
   );

  aliasv xaliasv79_ch8 (
    .PLUS(nd_aib79_ch2_x0y1),
    .MINUS(m1_ch2_aib[79])
   );

  aliasv xaliasv78_ch8 (
    .PLUS(nd_aib78_ch2_x0y1),
    .MINUS(m1_ch2_aib[78])
   );

  aliasv xaliasv77_ch8 (
    .PLUS(nd_aib77_ch2_x0y1),
    .MINUS(m1_ch2_aib[77])
   );

  aliasv xaliasv76_ch8 (
    .PLUS(nd_aib76_ch2_x0y1),
    .MINUS(m1_ch2_aib[76])
   );

  aliasv xaliasv75_ch8 (
    .PLUS(nd_aib75_ch2_x0y1),
    .MINUS(m1_ch2_aib[75])
   );

  aliasv xaliasv74_ch8 (
    .PLUS(nd_aib74_ch2_x0y1),
    .MINUS(m1_ch2_aib[74])
   );

  aliasv xaliasv73_ch8 (
    .PLUS(nd_aib73_ch2_x0y1),
    .MINUS(m1_ch2_aib[73])
   );

  aliasv xaliasv72_ch8 (
    .PLUS(nd_aib72_ch2_x0y1),
    .MINUS(m1_ch2_aib[72])
   );

  aliasv xaliasv71_ch8 (
    .PLUS(nd_aib71_ch2_x0y1),
    .MINUS(m1_ch2_aib[71])
   );

  aliasv xaliasv70_ch8 (
    .PLUS(nd_aib70_ch2_x0y1),
    .MINUS(m1_ch2_aib[70])
   );

  aliasv xaliasv69_ch8 (
    .PLUS(nd_aib69_ch2_x0y1),
    .MINUS(m1_ch2_aib[69])
   );

  aliasv xaliasv68_ch8 (
    .PLUS(nd_aib68_ch2_x0y1),
    .MINUS(m1_ch2_aib[68])
   );

  aliasv xaliasv67_ch8 (
    .PLUS(nd_aib67_ch2_x0y1),
    .MINUS(m1_ch2_aib[67])
   );

  aliasv xaliasv66_ch8 (
    .PLUS(nd_aib66_ch2_x0y1),
    .MINUS(m1_ch2_aib[66])
   );

  aliasv xaliasv65_ch8 (
    .PLUS(nd_aib65_ch2_x0y1),
    .MINUS(m1_ch2_aib[65])
   );

  aliasv xaliasv64_ch8 (
    .PLUS(nd_aib64_ch2_x0y1),
    .MINUS(m1_ch2_aib[64])
   );

  aliasv xaliasv63_ch8 (
    .PLUS(nd_aib63_ch2_x0y1),
    .MINUS(m1_ch2_aib[63])
   );

  aliasv xaliasv62_ch8 (
    .PLUS(nd_aib62_ch2_x0y1),
    .MINUS(m1_ch2_aib[62])
   );

  aliasv xaliasv61_ch8 (
    .PLUS(nd_aib61_ch2_x0y1),
    .MINUS(m1_ch2_aib[61])
   );

  aliasv xaliasv60_ch8 (
    .PLUS(nd_aib60_ch2_x0y1),
    .MINUS(m1_ch2_aib[60])
   );

  aliasv xaliasv59_ch8 (
    .PLUS(nd_aib59_ch2_x0y1),
    .MINUS(m1_ch2_aib[59])
   );

  aliasv xaliasv58_ch8 (
    .PLUS(nd_aib58_ch2_x0y1),
    .MINUS(m1_ch2_aib[58])
   );

  aliasv xaliasv57_ch8 (
    .PLUS(nd_aib57_ch2_x0y1),
    .MINUS(m1_ch2_aib[57])
   );

  aliasv xaliasv56_ch8 (
    .PLUS(nd_aib56_ch2_x0y1),
    .MINUS(m1_ch2_aib[56])
   );

  aliasv xaliasv55_ch8 (
    .PLUS(nd_aib55_ch2_x0y1),
    .MINUS(m1_ch2_aib[55])
   );

  aliasv xaliasv54_ch8 (
    .PLUS(nd_aib54_ch2_x0y1),
    .MINUS(m1_ch2_aib[54])
   );

  aliasv xaliasv53_ch8 (
    .PLUS(nd_aib53_ch2_x0y1),
    .MINUS(m1_ch2_aib[53])
   );

  aliasv xaliasv52_ch8 (
    .PLUS(nd_aib52_ch2_x0y1),
    .MINUS(m1_ch2_aib[52])
   );

  aliasv xaliasv51_ch8 (
    .PLUS(nd_aib51_ch2_x0y1),
    .MINUS(m1_ch2_aib[51])
   );

  aliasv xaliasv50_ch8 (
    .PLUS(nd_aib50_ch2_x0y1),
    .MINUS(m1_ch2_aib[50])
   );

  aliasv xaliasv49_ch8 (
    .PLUS(nd_aib49_ch2_x0y1),
    .MINUS(m1_ch2_aib[49])
   );

  aliasv xaliasv48_ch8 (
    .PLUS(nd_aib48_ch2_x0y1),
    .MINUS(m1_ch2_aib[48])
   );

  aliasv xaliasv47_ch8 (
    .PLUS(nd_aib47_ch2_x0y1),
    .MINUS(m1_ch2_aib[47])
   );

  aliasv xaliasv46_ch8 (
    .PLUS(nd_aib46_ch2_x0y1),
    .MINUS(m1_ch2_aib[46])
   );

  aliasv xaliasv45_ch8 (
    .PLUS(nd_aib45_ch2_x0y1),
    .MINUS(m1_ch2_aib[45])
   );

  aliasv xaliasv44_ch8 (
    .PLUS(nd_aib44_ch2_x0y1),
    .MINUS(m1_ch2_aib[44])
   );

  aliasv xaliasv43_ch8 (
    .PLUS(nd_aib43_ch2_x0y1),
    .MINUS(m1_ch2_aib[43])
   );

  aliasv xaliasv42_ch8 (
    .PLUS(nd_aib42_ch2_x0y1),
    .MINUS(m1_ch2_aib[42])
   );

  aliasv xaliasv41_ch8 (
    .PLUS(nd_aib41_ch2_x0y1),
    .MINUS(m1_ch2_aib[41])
   );

  aliasv xaliasv40_ch8 (
    .PLUS(nd_aib40_ch2_x0y1),
    .MINUS(m1_ch2_aib[40])
   );

  aliasv xaliasv39_ch8 (
    .PLUS(nd_aib39_ch2_x0y1),
    .MINUS(m1_ch2_aib[39])
   );

  aliasv xaliasv38_ch8 (
    .PLUS(nd_aib38_ch2_x0y1),
    .MINUS(m1_ch2_aib[38])
   );

  aliasv xaliasv37_ch8 (
    .PLUS(nd_aib37_ch2_x0y1),
    .MINUS(m1_ch2_aib[37])
   );

  aliasv xaliasv36_ch8 (
    .PLUS(nd_aib36_ch2_x0y1),
    .MINUS(m1_ch2_aib[36])
   );

  aliasv xaliasv35_ch8 (
    .PLUS(nd_aib35_ch2_x0y1),
    .MINUS(m1_ch2_aib[35])
   );

  aliasv xaliasv34_ch8 (
    .PLUS(nd_aib34_ch2_x0y1),
    .MINUS(m1_ch2_aib[34])
   );

  aliasv xaliasv33_ch8 (
    .PLUS(nd_aib33_ch2_x0y1),
    .MINUS(m1_ch2_aib[33])
   );

  aliasv xaliasv32_ch8 (
    .PLUS(nd_aib32_ch2_x0y1),
    .MINUS(m1_ch2_aib[32])
   );

  aliasv xaliasv31_ch8 (
    .PLUS(nd_aib31_ch2_x0y1),
    .MINUS(m1_ch2_aib[31])
   );

  aliasv xaliasv30_ch8 (
    .PLUS(nd_aib30_ch2_x0y1),
    .MINUS(m1_ch2_aib[30])
   );

  aliasv xaliasv29_ch8 (
    .PLUS(nd_aib29_ch2_x0y1),
    .MINUS(m1_ch2_aib[29])
   );

  aliasv xaliasv28_ch8 (
    .PLUS(nd_aib28_ch2_x0y1),
    .MINUS(m1_ch2_aib[28])
   );

  aliasv xaliasv27_ch8 (
    .PLUS(nd_aib27_ch2_x0y1),
    .MINUS(m1_ch2_aib[27])
   );

  aliasv xaliasv26_ch8 (
    .PLUS(nd_aib26_ch2_x0y1),
    .MINUS(m1_ch2_aib[26])
   );

  aliasv xaliasv25_ch8 (
    .PLUS(nd_aib25_ch2_x0y1),
    .MINUS(m1_ch2_aib[25])
   );

  aliasv xaliasv24_ch8 (
    .PLUS(nd_aib24_ch2_x0y1),
    .MINUS(m1_ch2_aib[24])
   );

  aliasv xaliasv23_ch8 (
    .PLUS(nd_aib23_ch2_x0y1),
    .MINUS(m1_ch2_aib[23])
   );

  aliasv xaliasv22_ch8 (
    .PLUS(nd_aib22_ch2_x0y1),
    .MINUS(m1_ch2_aib[22])
   );

  aliasv xaliasv21_ch8 (
    .PLUS(nd_aib21_ch2_x0y1),
    .MINUS(m1_ch2_aib[21])
   );

  aliasv xaliasv20_ch8 (
    .PLUS(nd_aib20_ch2_x0y1),
    .MINUS(m1_ch2_aib[20])
   );

  aliasv xaliasv19_ch8 (
    .PLUS(nd_aib19_ch2_x0y1),
    .MINUS(m1_ch2_aib[19])
   );

  aliasv xaliasv18_ch8 (
    .PLUS(nd_aib18_ch2_x0y1),
    .MINUS(m1_ch2_aib[18])
   );

  aliasv xaliasv17_ch8 (
    .PLUS(nd_aib17_ch2_x0y1),
    .MINUS(m1_ch2_aib[17])
   );

  aliasv xaliasv16_ch8 (
    .PLUS(nd_aib16_ch2_x0y1),
    .MINUS(m1_ch2_aib[16])
   );

  aliasv xaliasv15_ch8 (
    .PLUS(nd_aib15_ch2_x0y1),
    .MINUS(m1_ch2_aib[15])
   );

  aliasv xaliasv14_ch8 (
    .PLUS(nd_aib14_ch2_x0y1),
    .MINUS(m1_ch2_aib[14])
   );

  aliasv xaliasv13_ch8 (
    .PLUS(nd_aib13_ch2_x0y1),
    .MINUS(m1_ch2_aib[13])
   );

  aliasv xaliasv12_ch8 (
    .PLUS(nd_aib12_ch2_x0y1),
    .MINUS(m1_ch2_aib[12])
   );

  aliasv xaliasv11_ch8 (
    .PLUS(nd_aib11_ch2_x0y1),
    .MINUS(m1_ch2_aib[11])
   );

  aliasv xaliasv10_ch8 (
    .PLUS(nd_aib10_ch2_x0y1),
    .MINUS(m1_ch2_aib[10])
   );

  aliasv xaliasv9_ch8 (
    .PLUS(nd_aib9_ch2_x0y1),
    .MINUS(m1_ch2_aib[9])
   );

  aliasv xaliasv8_ch8 (
    .PLUS(nd_aib8_ch2_x0y1),
    .MINUS(m1_ch2_aib[8])
   );

  aliasv xaliasv7_ch8 (
    .PLUS(nd_aib7_ch2_x0y1),
    .MINUS(m1_ch2_aib[7])
   );

  aliasv xaliasv6_ch8 (
    .PLUS(nd_aib6_ch2_x0y1),
    .MINUS(m1_ch2_aib[6])
   );

  aliasv xaliasv5_ch8 (
    .PLUS(nd_aib5_ch2_x0y1),
    .MINUS(m1_ch2_aib[5])
   );

  aliasv xaliasv4_ch8 (
    .PLUS(nd_aib4_ch2_x0y1),
    .MINUS(m1_ch2_aib[4])
   );

  aliasv xaliasv3_ch8 (
    .PLUS(nd_aib3_ch2_x0y1),
    .MINUS(m1_ch2_aib[3])
   );

  aliasv xaliasv2_ch8 (
    .PLUS(nd_aib2_ch2_x0y1),
    .MINUS(m1_ch2_aib[2])
   );

  aliasv xaliasv1_ch8 (
    .PLUS(nd_aib1_ch2_x0y1),
    .MINUS(m1_ch2_aib[1])
   );

  aliasv xaliasv0_ch8 (
    .PLUS(nd_aib0_ch2_x0y1),
    .MINUS(m1_ch2_aib[0])
   );

// ## START OF  ch9 ( ##
  aliasv xaliasv95_ch9 (
    .PLUS(nd_aib95_ch3_x0y1),
    .MINUS(m1_ch3_aib[95])
   );

  aliasv xaliasv94_ch9 (
    .PLUS(nd_aib94_ch3_x0y1),
    .MINUS(m1_ch3_aib[94])
   );

  aliasv xaliasv93_ch9 (
    .PLUS(nd_aib93_ch3_x0y1),
    .MINUS(m1_ch3_aib[93])
   );

  aliasv xaliasv92_ch9 (
    .PLUS(nd_aib92_ch3_x0y1),
    .MINUS(m1_ch3_aib[92])
   );

  aliasv xaliasv91_ch9 (
    .PLUS(nd_aib91_ch3_x0y1),
    .MINUS(m1_ch3_aib[91])
   );

  aliasv xaliasv90_ch9 (
    .PLUS(nd_aib90_ch3_x0y1),
    .MINUS(m1_ch3_aib[90])
   );

  aliasv xaliasv89_ch9 (
    .PLUS(nd_aib89_ch3_x0y1),
    .MINUS(m1_ch3_aib[89])
   );

  aliasv xaliasv88_ch9 (
    .PLUS(nd_aib88_ch3_x0y1),
    .MINUS(m1_ch3_aib[88])
   );

  aliasv xaliasv87_ch9 (
    .PLUS(nd_aib87_ch3_x0y1),
    .MINUS(m1_ch3_aib[87])
   );

  aliasv xaliasv86_ch9 (
    .PLUS(nd_aib86_ch3_x0y1),
    .MINUS(m1_ch3_aib[86])
   );

  aliasv xaliasv85_ch9 (
    .PLUS(nd_aib85_ch3_x0y1),
    .MINUS(m1_ch3_aib[85])
   );

  aliasv xaliasv84_ch9 (
    .PLUS(nd_aib84_ch3_x0y1),
    .MINUS(m1_ch3_aib[84])
   );

  aliasv xaliasv83_ch9 (
    .PLUS(nd_aib83_ch3_x0y1),
    .MINUS(m1_ch3_aib[83])
   );

  aliasv xaliasv82_ch9 (
    .PLUS(nd_aib82_ch3_x0y1),
    .MINUS(m1_ch3_aib[82])
   );

  aliasv xaliasv81_ch9 (
    .PLUS(nd_aib81_ch3_x0y1),
    .MINUS(m1_ch3_aib[81])
   );

  aliasv xaliasv80_ch9 (
    .PLUS(nd_aib80_ch3_x0y1),
    .MINUS(m1_ch3_aib[80])
   );

  aliasv xaliasv79_ch9 (
    .PLUS(nd_aib79_ch3_x0y1),
    .MINUS(m1_ch3_aib[79])
   );

  aliasv xaliasv78_ch9 (
    .PLUS(nd_aib78_ch3_x0y1),
    .MINUS(m1_ch3_aib[78])
   );

  aliasv xaliasv77_ch9 (
    .PLUS(nd_aib77_ch3_x0y1),
    .MINUS(m1_ch3_aib[77])
   );

  aliasv xaliasv76_ch9 (
    .PLUS(nd_aib76_ch3_x0y1),
    .MINUS(m1_ch3_aib[76])
   );

  aliasv xaliasv75_ch9 (
    .PLUS(nd_aib75_ch3_x0y1),
    .MINUS(m1_ch3_aib[75])
   );

  aliasv xaliasv74_ch9 (
    .PLUS(nd_aib74_ch3_x0y1),
    .MINUS(m1_ch3_aib[74])
   );

  aliasv xaliasv73_ch9 (
    .PLUS(nd_aib73_ch3_x0y1),
    .MINUS(m1_ch3_aib[73])
   );

  aliasv xaliasv72_ch9 (
    .PLUS(nd_aib72_ch3_x0y1),
    .MINUS(m1_ch3_aib[72])
   );

  aliasv xaliasv71_ch9 (
    .PLUS(nd_aib71_ch3_x0y1),
    .MINUS(m1_ch3_aib[71])
   );

  aliasv xaliasv70_ch9 (
    .PLUS(nd_aib70_ch3_x0y1),
    .MINUS(m1_ch3_aib[70])
   );

  aliasv xaliasv69_ch9 (
    .PLUS(nd_aib69_ch3_x0y1),
    .MINUS(m1_ch3_aib[69])
   );

  aliasv xaliasv68_ch9 (
    .PLUS(nd_aib68_ch3_x0y1),
    .MINUS(m1_ch3_aib[68])
   );

  aliasv xaliasv67_ch9 (
    .PLUS(nd_aib67_ch3_x0y1),
    .MINUS(m1_ch3_aib[67])
   );

  aliasv xaliasv66_ch9 (
    .PLUS(nd_aib66_ch3_x0y1),
    .MINUS(m1_ch3_aib[66])
   );

  aliasv xaliasv65_ch9 (
    .PLUS(nd_aib65_ch3_x0y1),
    .MINUS(m1_ch3_aib[65])
   );

  aliasv xaliasv64_ch9 (
    .PLUS(nd_aib64_ch3_x0y1),
    .MINUS(m1_ch3_aib[64])
   );

  aliasv xaliasv63_ch9 (
    .PLUS(nd_aib63_ch3_x0y1),
    .MINUS(m1_ch3_aib[63])
   );

  aliasv xaliasv62_ch9 (
    .PLUS(nd_aib62_ch3_x0y1),
    .MINUS(m1_ch3_aib[62])
   );

  aliasv xaliasv61_ch9 (
    .PLUS(nd_aib61_ch3_x0y1),
    .MINUS(m1_ch3_aib[61])
   );

  aliasv xaliasv60_ch9 (
    .PLUS(nd_aib60_ch3_x0y1),
    .MINUS(m1_ch3_aib[60])
   );

  aliasv xaliasv59_ch9 (
    .PLUS(nd_aib59_ch3_x0y1),
    .MINUS(m1_ch3_aib[59])
   );

  aliasv xaliasv58_ch9 (
    .PLUS(nd_aib58_ch3_x0y1),
    .MINUS(m1_ch3_aib[58])
   );

  aliasv xaliasv57_ch9 (
    .PLUS(nd_aib57_ch3_x0y1),
    .MINUS(m1_ch3_aib[57])
   );

  aliasv xaliasv56_ch9 (
    .PLUS(nd_aib56_ch3_x0y1),
    .MINUS(m1_ch3_aib[56])
   );

  aliasv xaliasv55_ch9 (
    .PLUS(nd_aib55_ch3_x0y1),
    .MINUS(m1_ch3_aib[55])
   );

  aliasv xaliasv54_ch9 (
    .PLUS(nd_aib54_ch3_x0y1),
    .MINUS(m1_ch3_aib[54])
   );

  aliasv xaliasv53_ch9 (
    .PLUS(nd_aib53_ch3_x0y1),
    .MINUS(m1_ch3_aib[53])
   );

  aliasv xaliasv52_ch9 (
    .PLUS(nd_aib52_ch3_x0y1),
    .MINUS(m1_ch3_aib[52])
   );

  aliasv xaliasv51_ch9 (
    .PLUS(nd_aib51_ch3_x0y1),
    .MINUS(m1_ch3_aib[51])
   );

  aliasv xaliasv50_ch9 (
    .PLUS(nd_aib50_ch3_x0y1),
    .MINUS(m1_ch3_aib[50])
   );

  aliasv xaliasv49_ch9 (
    .PLUS(nd_aib49_ch3_x0y1),
    .MINUS(m1_ch3_aib[49])
   );

  aliasv xaliasv48_ch9 (
    .PLUS(nd_aib48_ch3_x0y1),
    .MINUS(m1_ch3_aib[48])
   );

  aliasv xaliasv47_ch9 (
    .PLUS(nd_aib47_ch3_x0y1),
    .MINUS(m1_ch3_aib[47])
   );

  aliasv xaliasv46_ch9 (
    .PLUS(nd_aib46_ch3_x0y1),
    .MINUS(m1_ch3_aib[46])
   );

  aliasv xaliasv45_ch9 (
    .PLUS(nd_aib45_ch3_x0y1),
    .MINUS(m1_ch3_aib[45])
   );

  aliasv xaliasv44_ch9 (
    .PLUS(nd_aib44_ch3_x0y1),
    .MINUS(m1_ch3_aib[44])
   );

  aliasv xaliasv43_ch9 (
    .PLUS(nd_aib43_ch3_x0y1),
    .MINUS(m1_ch3_aib[43])
   );

  aliasv xaliasv42_ch9 (
    .PLUS(nd_aib42_ch3_x0y1),
    .MINUS(m1_ch3_aib[42])
   );

  aliasv xaliasv41_ch9 (
    .PLUS(nd_aib41_ch3_x0y1),
    .MINUS(m1_ch3_aib[41])
   );

  aliasv xaliasv40_ch9 (
    .PLUS(nd_aib40_ch3_x0y1),
    .MINUS(m1_ch3_aib[40])
   );

  aliasv xaliasv39_ch9 (
    .PLUS(nd_aib39_ch3_x0y1),
    .MINUS(m1_ch3_aib[39])
   );

  aliasv xaliasv38_ch9 (
    .PLUS(nd_aib38_ch3_x0y1),
    .MINUS(m1_ch3_aib[38])
   );

  aliasv xaliasv37_ch9 (
    .PLUS(nd_aib37_ch3_x0y1),
    .MINUS(m1_ch3_aib[37])
   );

  aliasv xaliasv36_ch9 (
    .PLUS(nd_aib36_ch3_x0y1),
    .MINUS(m1_ch3_aib[36])
   );

  aliasv xaliasv35_ch9 (
    .PLUS(nd_aib35_ch3_x0y1),
    .MINUS(m1_ch3_aib[35])
   );

  aliasv xaliasv34_ch9 (
    .PLUS(nd_aib34_ch3_x0y1),
    .MINUS(m1_ch3_aib[34])
   );

  aliasv xaliasv33_ch9 (
    .PLUS(nd_aib33_ch3_x0y1),
    .MINUS(m1_ch3_aib[33])
   );

  aliasv xaliasv32_ch9 (
    .PLUS(nd_aib32_ch3_x0y1),
    .MINUS(m1_ch3_aib[32])
   );

  aliasv xaliasv31_ch9 (
    .PLUS(nd_aib31_ch3_x0y1),
    .MINUS(m1_ch3_aib[31])
   );

  aliasv xaliasv30_ch9 (
    .PLUS(nd_aib30_ch3_x0y1),
    .MINUS(m1_ch3_aib[30])
   );

  aliasv xaliasv29_ch9 (
    .PLUS(nd_aib29_ch3_x0y1),
    .MINUS(m1_ch3_aib[29])
   );

  aliasv xaliasv28_ch9 (
    .PLUS(nd_aib28_ch3_x0y1),
    .MINUS(m1_ch3_aib[28])
   );

  aliasv xaliasv27_ch9 (
    .PLUS(nd_aib27_ch3_x0y1),
    .MINUS(m1_ch3_aib[27])
   );

  aliasv xaliasv26_ch9 (
    .PLUS(nd_aib26_ch3_x0y1),
    .MINUS(m1_ch3_aib[26])
   );

  aliasv xaliasv25_ch9 (
    .PLUS(nd_aib25_ch3_x0y1),
    .MINUS(m1_ch3_aib[25])
   );

  aliasv xaliasv24_ch9 (
    .PLUS(nd_aib24_ch3_x0y1),
    .MINUS(m1_ch3_aib[24])
   );

  aliasv xaliasv23_ch9 (
    .PLUS(nd_aib23_ch3_x0y1),
    .MINUS(m1_ch3_aib[23])
   );

  aliasv xaliasv22_ch9 (
    .PLUS(nd_aib22_ch3_x0y1),
    .MINUS(m1_ch3_aib[22])
   );

  aliasv xaliasv21_ch9 (
    .PLUS(nd_aib21_ch3_x0y1),
    .MINUS(m1_ch3_aib[21])
   );

  aliasv xaliasv20_ch9 (
    .PLUS(nd_aib20_ch3_x0y1),
    .MINUS(m1_ch3_aib[20])
   );

  aliasv xaliasv19_ch9 (
    .PLUS(nd_aib19_ch3_x0y1),
    .MINUS(m1_ch3_aib[19])
   );

  aliasv xaliasv18_ch9 (
    .PLUS(nd_aib18_ch3_x0y1),
    .MINUS(m1_ch3_aib[18])
   );

  aliasv xaliasv17_ch9 (
    .PLUS(nd_aib17_ch3_x0y1),
    .MINUS(m1_ch3_aib[17])
   );

  aliasv xaliasv16_ch9 (
    .PLUS(nd_aib16_ch3_x0y1),
    .MINUS(m1_ch3_aib[16])
   );

  aliasv xaliasv15_ch9 (
    .PLUS(nd_aib15_ch3_x0y1),
    .MINUS(m1_ch3_aib[15])
   );

  aliasv xaliasv14_ch9 (
    .PLUS(nd_aib14_ch3_x0y1),
    .MINUS(m1_ch3_aib[14])
   );

  aliasv xaliasv13_ch9 (
    .PLUS(nd_aib13_ch3_x0y1),
    .MINUS(m1_ch3_aib[13])
   );

  aliasv xaliasv12_ch9 (
    .PLUS(nd_aib12_ch3_x0y1),
    .MINUS(m1_ch3_aib[12])
   );

  aliasv xaliasv11_ch9 (
    .PLUS(nd_aib11_ch3_x0y1),
    .MINUS(m1_ch3_aib[11])
   );

  aliasv xaliasv10_ch9 (
    .PLUS(nd_aib10_ch3_x0y1),
    .MINUS(m1_ch3_aib[10])
   );

  aliasv xaliasv9_ch9 (
    .PLUS(nd_aib9_ch3_x0y1),
    .MINUS(m1_ch3_aib[9])
   );

  aliasv xaliasv8_ch9 (
    .PLUS(nd_aib8_ch3_x0y1),
    .MINUS(m1_ch3_aib[8])
   );

  aliasv xaliasv7_ch9 (
    .PLUS(nd_aib7_ch3_x0y1),
    .MINUS(m1_ch3_aib[7])
   );

  aliasv xaliasv6_ch9 (
    .PLUS(nd_aib6_ch3_x0y1),
    .MINUS(m1_ch3_aib[6])
   );

  aliasv xaliasv5_ch9 (
    .PLUS(nd_aib5_ch3_x0y1),
    .MINUS(m1_ch3_aib[5])
   );

  aliasv xaliasv4_ch9 (
    .PLUS(nd_aib4_ch3_x0y1),
    .MINUS(m1_ch3_aib[4])
   );

  aliasv xaliasv3_ch9 (
    .PLUS(nd_aib3_ch3_x0y1),
    .MINUS(m1_ch3_aib[3])
   );

  aliasv xaliasv2_ch9 (
    .PLUS(nd_aib2_ch3_x0y1),
    .MINUS(m1_ch3_aib[2])
   );

  aliasv xaliasv1_ch9 (
    .PLUS(nd_aib1_ch3_x0y1),
    .MINUS(m1_ch3_aib[1])
   );

  aliasv xaliasv0_ch9 (
    .PLUS(nd_aib0_ch3_x0y1),
    .MINUS(m1_ch3_aib[0])
   );

// ## START OF  ch10 ( ##
  aliasv xaliasv95_ch10 (
    .PLUS(nd_aib95_ch4_x0y1),
    .MINUS(m1_ch4_aib[95])
   );

  aliasv xaliasv94_ch10 (
    .PLUS(nd_aib94_ch4_x0y1),
    .MINUS(m1_ch4_aib[94])
   );

  aliasv xaliasv93_ch10 (
    .PLUS(nd_aib93_ch4_x0y1),
    .MINUS(m1_ch4_aib[93])
   );

  aliasv xaliasv92_ch10 (
    .PLUS(nd_aib92_ch4_x0y1),
    .MINUS(m1_ch4_aib[92])
   );

  aliasv xaliasv91_ch10 (
    .PLUS(nd_aib91_ch4_x0y1),
    .MINUS(m1_ch4_aib[91])
   );

  aliasv xaliasv90_ch10 (
    .PLUS(nd_aib90_ch4_x0y1),
    .MINUS(m1_ch4_aib[90])
   );

  aliasv xaliasv89_ch10 (
    .PLUS(nd_aib89_ch4_x0y1),
    .MINUS(m1_ch4_aib[89])
   );

  aliasv xaliasv88_ch10 (
    .PLUS(nd_aib88_ch4_x0y1),
    .MINUS(m1_ch4_aib[88])
   );

  aliasv xaliasv87_ch10 (
    .PLUS(nd_aib87_ch4_x0y1),
    .MINUS(m1_ch4_aib[87])
   );

  aliasv xaliasv86_ch10 (
    .PLUS(nd_aib86_ch4_x0y1),
    .MINUS(m1_ch4_aib[86])
   );

  aliasv xaliasv85_ch10 (
    .PLUS(nd_aib85_ch4_x0y1),
    .MINUS(m1_ch4_aib[85])
   );

  aliasv xaliasv84_ch10 (
    .PLUS(nd_aib84_ch4_x0y1),
    .MINUS(m1_ch4_aib[84])
   );

  aliasv xaliasv83_ch10 (
    .PLUS(nd_aib83_ch4_x0y1),
    .MINUS(m1_ch4_aib[83])
   );

  aliasv xaliasv82_ch10 (
    .PLUS(nd_aib82_ch4_x0y1),
    .MINUS(m1_ch4_aib[82])
   );

  aliasv xaliasv81_ch10 (
    .PLUS(nd_aib81_ch4_x0y1),
    .MINUS(m1_ch4_aib[81])
   );

  aliasv xaliasv80_ch10 (
    .PLUS(nd_aib80_ch4_x0y1),
    .MINUS(m1_ch4_aib[80])
   );

  aliasv xaliasv79_ch10 (
    .PLUS(nd_aib79_ch4_x0y1),
    .MINUS(m1_ch4_aib[79])
   );

  aliasv xaliasv78_ch10 (
    .PLUS(nd_aib78_ch4_x0y1),
    .MINUS(m1_ch4_aib[78])
   );

  aliasv xaliasv77_ch10 (
    .PLUS(nd_aib77_ch4_x0y1),
    .MINUS(m1_ch4_aib[77])
   );

  aliasv xaliasv76_ch10 (
    .PLUS(nd_aib76_ch4_x0y1),
    .MINUS(m1_ch4_aib[76])
   );

  aliasv xaliasv75_ch10 (
    .PLUS(nd_aib75_ch4_x0y1),
    .MINUS(m1_ch4_aib[75])
   );

  aliasv xaliasv74_ch10 (
    .PLUS(nd_aib74_ch4_x0y1),
    .MINUS(m1_ch4_aib[74])
   );

  aliasv xaliasv73_ch10 (
    .PLUS(nd_aib73_ch4_x0y1),
    .MINUS(m1_ch4_aib[73])
   );

  aliasv xaliasv72_ch10 (
    .PLUS(nd_aib72_ch4_x0y1),
    .MINUS(m1_ch4_aib[72])
   );

  aliasv xaliasv71_ch10 (
    .PLUS(nd_aib71_ch4_x0y1),
    .MINUS(m1_ch4_aib[71])
   );

  aliasv xaliasv70_ch10 (
    .PLUS(nd_aib70_ch4_x0y1),
    .MINUS(m1_ch4_aib[70])
   );

  aliasv xaliasv69_ch10 (
    .PLUS(nd_aib69_ch4_x0y1),
    .MINUS(m1_ch4_aib[69])
   );

  aliasv xaliasv68_ch10 (
    .PLUS(nd_aib68_ch4_x0y1),
    .MINUS(m1_ch4_aib[68])
   );

  aliasv xaliasv67_ch10 (
    .PLUS(nd_aib67_ch4_x0y1),
    .MINUS(m1_ch4_aib[67])
   );

  aliasv xaliasv66_ch10 (
    .PLUS(nd_aib66_ch4_x0y1),
    .MINUS(m1_ch4_aib[66])
   );

  aliasv xaliasv65_ch10 (
    .PLUS(nd_aib65_ch4_x0y1),
    .MINUS(m1_ch4_aib[65])
   );

  aliasv xaliasv64_ch10 (
    .PLUS(nd_aib64_ch4_x0y1),
    .MINUS(m1_ch4_aib[64])
   );

  aliasv xaliasv63_ch10 (
    .PLUS(nd_aib63_ch4_x0y1),
    .MINUS(m1_ch4_aib[63])
   );

  aliasv xaliasv62_ch10 (
    .PLUS(nd_aib62_ch4_x0y1),
    .MINUS(m1_ch4_aib[62])
   );

  aliasv xaliasv61_ch10 (
    .PLUS(nd_aib61_ch4_x0y1),
    .MINUS(m1_ch4_aib[61])
   );

  aliasv xaliasv60_ch10 (
    .PLUS(nd_aib60_ch4_x0y1),
    .MINUS(m1_ch4_aib[60])
   );

  aliasv xaliasv59_ch10 (
    .PLUS(nd_aib59_ch4_x0y1),
    .MINUS(m1_ch4_aib[59])
   );

  aliasv xaliasv58_ch10 (
    .PLUS(nd_aib58_ch4_x0y1),
    .MINUS(m1_ch4_aib[58])
   );

  aliasv xaliasv57_ch10 (
    .PLUS(nd_aib57_ch4_x0y1),
    .MINUS(m1_ch4_aib[57])
   );

  aliasv xaliasv56_ch10 (
    .PLUS(nd_aib56_ch4_x0y1),
    .MINUS(m1_ch4_aib[56])
   );

  aliasv xaliasv55_ch10 (
    .PLUS(nd_aib55_ch4_x0y1),
    .MINUS(m1_ch4_aib[55])
   );

  aliasv xaliasv54_ch10 (
    .PLUS(nd_aib54_ch4_x0y1),
    .MINUS(m1_ch4_aib[54])
   );

  aliasv xaliasv53_ch10 (
    .PLUS(nd_aib53_ch4_x0y1),
    .MINUS(m1_ch4_aib[53])
   );

  aliasv xaliasv52_ch10 (
    .PLUS(nd_aib52_ch4_x0y1),
    .MINUS(m1_ch4_aib[52])
   );

  aliasv xaliasv51_ch10 (
    .PLUS(nd_aib51_ch4_x0y1),
    .MINUS(m1_ch4_aib[51])
   );

  aliasv xaliasv50_ch10 (
    .PLUS(nd_aib50_ch4_x0y1),
    .MINUS(m1_ch4_aib[50])
   );

  aliasv xaliasv49_ch10 (
    .PLUS(nd_aib49_ch4_x0y1),
    .MINUS(m1_ch4_aib[49])
   );

  aliasv xaliasv48_ch10 (
    .PLUS(nd_aib48_ch4_x0y1),
    .MINUS(m1_ch4_aib[48])
   );

  aliasv xaliasv47_ch10 (
    .PLUS(nd_aib47_ch4_x0y1),
    .MINUS(m1_ch4_aib[47])
   );

  aliasv xaliasv46_ch10 (
    .PLUS(nd_aib46_ch4_x0y1),
    .MINUS(m1_ch4_aib[46])
   );

  aliasv xaliasv45_ch10 (
    .PLUS(nd_aib45_ch4_x0y1),
    .MINUS(m1_ch4_aib[45])
   );

  aliasv xaliasv44_ch10 (
    .PLUS(nd_aib44_ch4_x0y1),
    .MINUS(m1_ch4_aib[44])
   );

  aliasv xaliasv43_ch10 (
    .PLUS(nd_aib43_ch4_x0y1),
    .MINUS(m1_ch4_aib[43])
   );

  aliasv xaliasv42_ch10 (
    .PLUS(nd_aib42_ch4_x0y1),
    .MINUS(m1_ch4_aib[42])
   );

  aliasv xaliasv41_ch10 (
    .PLUS(nd_aib41_ch4_x0y1),
    .MINUS(m1_ch4_aib[41])
   );

  aliasv xaliasv40_ch10 (
    .PLUS(nd_aib40_ch4_x0y1),
    .MINUS(m1_ch4_aib[40])
   );

  aliasv xaliasv39_ch10 (
    .PLUS(nd_aib39_ch4_x0y1),
    .MINUS(m1_ch4_aib[39])
   );

  aliasv xaliasv38_ch10 (
    .PLUS(nd_aib38_ch4_x0y1),
    .MINUS(m1_ch4_aib[38])
   );

  aliasv xaliasv37_ch10 (
    .PLUS(nd_aib37_ch4_x0y1),
    .MINUS(m1_ch4_aib[37])
   );

  aliasv xaliasv36_ch10 (
    .PLUS(nd_aib36_ch4_x0y1),
    .MINUS(m1_ch4_aib[36])
   );

  aliasv xaliasv35_ch10 (
    .PLUS(nd_aib35_ch4_x0y1),
    .MINUS(m1_ch4_aib[35])
   );

  aliasv xaliasv34_ch10 (
    .PLUS(nd_aib34_ch4_x0y1),
    .MINUS(m1_ch4_aib[34])
   );

  aliasv xaliasv33_ch10 (
    .PLUS(nd_aib33_ch4_x0y1),
    .MINUS(m1_ch4_aib[33])
   );

  aliasv xaliasv32_ch10 (
    .PLUS(nd_aib32_ch4_x0y1),
    .MINUS(m1_ch4_aib[32])
   );

  aliasv xaliasv31_ch10 (
    .PLUS(nd_aib31_ch4_x0y1),
    .MINUS(m1_ch4_aib[31])
   );

  aliasv xaliasv30_ch10 (
    .PLUS(nd_aib30_ch4_x0y1),
    .MINUS(m1_ch4_aib[30])
   );

  aliasv xaliasv29_ch10 (
    .PLUS(nd_aib29_ch4_x0y1),
    .MINUS(m1_ch4_aib[29])
   );

  aliasv xaliasv28_ch10 (
    .PLUS(nd_aib28_ch4_x0y1),
    .MINUS(m1_ch4_aib[28])
   );

  aliasv xaliasv27_ch10 (
    .PLUS(nd_aib27_ch4_x0y1),
    .MINUS(m1_ch4_aib[27])
   );

  aliasv xaliasv26_ch10 (
    .PLUS(nd_aib26_ch4_x0y1),
    .MINUS(m1_ch4_aib[26])
   );

  aliasv xaliasv25_ch10 (
    .PLUS(nd_aib25_ch4_x0y1),
    .MINUS(m1_ch4_aib[25])
   );

  aliasv xaliasv24_ch10 (
    .PLUS(nd_aib24_ch4_x0y1),
    .MINUS(m1_ch4_aib[24])
   );

  aliasv xaliasv23_ch10 (
    .PLUS(nd_aib23_ch4_x0y1),
    .MINUS(m1_ch4_aib[23])
   );

  aliasv xaliasv22_ch10 (
    .PLUS(nd_aib22_ch4_x0y1),
    .MINUS(m1_ch4_aib[22])
   );

  aliasv xaliasv21_ch10 (
    .PLUS(nd_aib21_ch4_x0y1),
    .MINUS(m1_ch4_aib[21])
   );

  aliasv xaliasv20_ch10 (
    .PLUS(nd_aib20_ch4_x0y1),
    .MINUS(m1_ch4_aib[20])
   );

  aliasv xaliasv19_ch10 (
    .PLUS(nd_aib19_ch4_x0y1),
    .MINUS(m1_ch4_aib[19])
   );

  aliasv xaliasv18_ch10 (
    .PLUS(nd_aib18_ch4_x0y1),
    .MINUS(m1_ch4_aib[18])
   );

  aliasv xaliasv17_ch10 (
    .PLUS(nd_aib17_ch4_x0y1),
    .MINUS(m1_ch4_aib[17])
   );

  aliasv xaliasv16_ch10 (
    .PLUS(nd_aib16_ch4_x0y1),
    .MINUS(m1_ch4_aib[16])
   );

  aliasv xaliasv15_ch10 (
    .PLUS(nd_aib15_ch4_x0y1),
    .MINUS(m1_ch4_aib[15])
   );

  aliasv xaliasv14_ch10 (
    .PLUS(nd_aib14_ch4_x0y1),
    .MINUS(m1_ch4_aib[14])
   );

  aliasv xaliasv13_ch10 (
    .PLUS(nd_aib13_ch4_x0y1),
    .MINUS(m1_ch4_aib[13])
   );

  aliasv xaliasv12_ch10 (
    .PLUS(nd_aib12_ch4_x0y1),
    .MINUS(m1_ch4_aib[12])
   );

  aliasv xaliasv11_ch10 (
    .PLUS(nd_aib11_ch4_x0y1),
    .MINUS(m1_ch4_aib[11])
   );

  aliasv xaliasv10_ch10 (
    .PLUS(nd_aib10_ch4_x0y1),
    .MINUS(m1_ch4_aib[10])
   );

  aliasv xaliasv9_ch10 (
    .PLUS(nd_aib9_ch4_x0y1),
    .MINUS(m1_ch4_aib[9])
   );

  aliasv xaliasv8_ch10 (
    .PLUS(nd_aib8_ch4_x0y1),
    .MINUS(m1_ch4_aib[8])
   );

  aliasv xaliasv7_ch10 (
    .PLUS(nd_aib7_ch4_x0y1),
    .MINUS(m1_ch4_aib[7])
   );

  aliasv xaliasv6_ch10 (
    .PLUS(nd_aib6_ch4_x0y1),
    .MINUS(m1_ch4_aib[6])
   );

  aliasv xaliasv5_ch10 (
    .PLUS(nd_aib5_ch4_x0y1),
    .MINUS(m1_ch4_aib[5])
   );

  aliasv xaliasv4_ch10 (
    .PLUS(nd_aib4_ch4_x0y1),
    .MINUS(m1_ch4_aib[4])
   );

  aliasv xaliasv3_ch10 (
    .PLUS(nd_aib3_ch4_x0y1),
    .MINUS(m1_ch4_aib[3])
   );

  aliasv xaliasv2_ch10 (
    .PLUS(nd_aib2_ch4_x0y1),
    .MINUS(m1_ch4_aib[2])
   );

  aliasv xaliasv1_ch10 (
    .PLUS(nd_aib1_ch4_x0y1),
    .MINUS(m1_ch4_aib[1])
   );

  aliasv xaliasv0_ch10 (
    .PLUS(nd_aib0_ch4_x0y1),
    .MINUS(m1_ch4_aib[0])
   );

// ## START OF  ch11 ( ##
  aliasv xaliasv95_ch11 (
    .PLUS(nd_aib95_ch5_x0y1),
    .MINUS(m1_ch5_aib[95])
   );

  aliasv xaliasv94_ch11 (
    .PLUS(nd_aib94_ch5_x0y1),
    .MINUS(m1_ch5_aib[94])
   );

  aliasv xaliasv93_ch11 (
    .PLUS(nd_aib93_ch5_x0y1),
    .MINUS(m1_ch5_aib[93])
   );

  aliasv xaliasv92_ch11 (
    .PLUS(nd_aib92_ch5_x0y1),
    .MINUS(m1_ch5_aib[92])
   );

  aliasv xaliasv91_ch11 (
    .PLUS(nd_aib91_ch5_x0y1),
    .MINUS(m1_ch5_aib[91])
   );

  aliasv xaliasv90_ch11 (
    .PLUS(nd_aib90_ch5_x0y1),
    .MINUS(m1_ch5_aib[90])
   );

  aliasv xaliasv89_ch11 (
    .PLUS(nd_aib89_ch5_x0y1),
    .MINUS(m1_ch5_aib[89])
   );

  aliasv xaliasv88_ch11 (
    .PLUS(nd_aib88_ch5_x0y1),
    .MINUS(m1_ch5_aib[88])
   );

  aliasv xaliasv87_ch11 (
    .PLUS(nd_aib87_ch5_x0y1),
    .MINUS(m1_ch5_aib[87])
   );

  aliasv xaliasv86_ch11 (
    .PLUS(nd_aib86_ch5_x0y1),
    .MINUS(m1_ch5_aib[86])
   );

  aliasv xaliasv85_ch11 (
    .PLUS(nd_aib85_ch5_x0y1),
    .MINUS(m1_ch5_aib[85])
   );

  aliasv xaliasv84_ch11 (
    .PLUS(nd_aib84_ch5_x0y1),
    .MINUS(m1_ch5_aib[84])
   );

  aliasv xaliasv83_ch11 (
    .PLUS(nd_aib83_ch5_x0y1),
    .MINUS(m1_ch5_aib[83])
   );

  aliasv xaliasv82_ch11 (
    .PLUS(nd_aib82_ch5_x0y1),
    .MINUS(m1_ch5_aib[82])
   );

  aliasv xaliasv81_ch11 (
    .PLUS(nd_aib81_ch5_x0y1),
    .MINUS(m1_ch5_aib[81])
   );

  aliasv xaliasv80_ch11 (
    .PLUS(nd_aib80_ch5_x0y1),
    .MINUS(m1_ch5_aib[80])
   );

  aliasv xaliasv79_ch11 (
    .PLUS(nd_aib79_ch5_x0y1),
    .MINUS(m1_ch5_aib[79])
   );

  aliasv xaliasv78_ch11 (
    .PLUS(nd_aib78_ch5_x0y1),
    .MINUS(m1_ch5_aib[78])
   );

  aliasv xaliasv77_ch11 (
    .PLUS(nd_aib77_ch5_x0y1),
    .MINUS(m1_ch5_aib[77])
   );

  aliasv xaliasv76_ch11 (
    .PLUS(nd_aib76_ch5_x0y1),
    .MINUS(m1_ch5_aib[76])
   );

  aliasv xaliasv75_ch11 (
    .PLUS(nd_aib75_ch5_x0y1),
    .MINUS(m1_ch5_aib[75])
   );

  aliasv xaliasv74_ch11 (
    .PLUS(nd_aib74_ch5_x0y1),
    .MINUS(m1_ch5_aib[74])
   );

  aliasv xaliasv73_ch11 (
    .PLUS(nd_aib73_ch5_x0y1),
    .MINUS(m1_ch5_aib[73])
   );

  aliasv xaliasv72_ch11 (
    .PLUS(nd_aib72_ch5_x0y1),
    .MINUS(m1_ch5_aib[72])
   );

  aliasv xaliasv71_ch11 (
    .PLUS(nd_aib71_ch5_x0y1),
    .MINUS(m1_ch5_aib[71])
   );

  aliasv xaliasv70_ch11 (
    .PLUS(nd_aib70_ch5_x0y1),
    .MINUS(m1_ch5_aib[70])
   );

  aliasv xaliasv69_ch11 (
    .PLUS(nd_aib69_ch5_x0y1),
    .MINUS(m1_ch5_aib[69])
   );

  aliasv xaliasv68_ch11 (
    .PLUS(nd_aib68_ch5_x0y1),
    .MINUS(m1_ch5_aib[68])
   );

  aliasv xaliasv67_ch11 (
    .PLUS(nd_aib67_ch5_x0y1),
    .MINUS(m1_ch5_aib[67])
   );

  aliasv xaliasv66_ch11 (
    .PLUS(nd_aib66_ch5_x0y1),
    .MINUS(m1_ch5_aib[66])
   );

  aliasv xaliasv65_ch11 (
    .PLUS(nd_aib65_ch5_x0y1),
    .MINUS(m1_ch5_aib[65])
   );

  aliasv xaliasv64_ch11 (
    .PLUS(nd_aib64_ch5_x0y1),
    .MINUS(m1_ch5_aib[64])
   );

  aliasv xaliasv63_ch11 (
    .PLUS(nd_aib63_ch5_x0y1),
    .MINUS(m1_ch5_aib[63])
   );

  aliasv xaliasv62_ch11 (
    .PLUS(nd_aib62_ch5_x0y1),
    .MINUS(m1_ch5_aib[62])
   );

  aliasv xaliasv61_ch11 (
    .PLUS(nd_aib61_ch5_x0y1),
    .MINUS(m1_ch5_aib[61])
   );

  aliasv xaliasv60_ch11 (
    .PLUS(nd_aib60_ch5_x0y1),
    .MINUS(m1_ch5_aib[60])
   );

  aliasv xaliasv59_ch11 (
    .PLUS(nd_aib59_ch5_x0y1),
    .MINUS(m1_ch5_aib[59])
   );

  aliasv xaliasv58_ch11 (
    .PLUS(nd_aib58_ch5_x0y1),
    .MINUS(m1_ch5_aib[58])
   );

  aliasv xaliasv57_ch11 (
    .PLUS(nd_aib57_ch5_x0y1),
    .MINUS(m1_ch5_aib[57])
   );

  aliasv xaliasv56_ch11 (
    .PLUS(nd_aib56_ch5_x0y1),
    .MINUS(m1_ch5_aib[56])
   );

  aliasv xaliasv55_ch11 (
    .PLUS(nd_aib55_ch5_x0y1),
    .MINUS(m1_ch5_aib[55])
   );

  aliasv xaliasv54_ch11 (
    .PLUS(nd_aib54_ch5_x0y1),
    .MINUS(m1_ch5_aib[54])
   );

  aliasv xaliasv53_ch11 (
    .PLUS(nd_aib53_ch5_x0y1),
    .MINUS(m1_ch5_aib[53])
   );

  aliasv xaliasv52_ch11 (
    .PLUS(nd_aib52_ch5_x0y1),
    .MINUS(m1_ch5_aib[52])
   );

  aliasv xaliasv51_ch11 (
    .PLUS(nd_aib51_ch5_x0y1),
    .MINUS(m1_ch5_aib[51])
   );

  aliasv xaliasv50_ch11 (
    .PLUS(nd_aib50_ch5_x0y1),
    .MINUS(m1_ch5_aib[50])
   );

  aliasv xaliasv49_ch11 (
    .PLUS(nd_aib49_ch5_x0y1),
    .MINUS(m1_ch5_aib[49])
   );

  aliasv xaliasv48_ch11 (
    .PLUS(nd_aib48_ch5_x0y1),
    .MINUS(m1_ch5_aib[48])
   );

  aliasv xaliasv47_ch11 (
    .PLUS(nd_aib47_ch5_x0y1),
    .MINUS(m1_ch5_aib[47])
   );

  aliasv xaliasv46_ch11 (
    .PLUS(nd_aib46_ch5_x0y1),
    .MINUS(m1_ch5_aib[46])
   );

  aliasv xaliasv45_ch11 (
    .PLUS(nd_aib45_ch5_x0y1),
    .MINUS(m1_ch5_aib[45])
   );

  aliasv xaliasv44_ch11 (
    .PLUS(nd_aib44_ch5_x0y1),
    .MINUS(m1_ch5_aib[44])
   );

  aliasv xaliasv43_ch11 (
    .PLUS(nd_aib43_ch5_x0y1),
    .MINUS(m1_ch5_aib[43])
   );

  aliasv xaliasv42_ch11 (
    .PLUS(nd_aib42_ch5_x0y1),
    .MINUS(m1_ch5_aib[42])
   );

  aliasv xaliasv41_ch11 (
    .PLUS(nd_aib41_ch5_x0y1),
    .MINUS(m1_ch5_aib[41])
   );

  aliasv xaliasv40_ch11 (
    .PLUS(nd_aib40_ch5_x0y1),
    .MINUS(m1_ch5_aib[40])
   );

  aliasv xaliasv39_ch11 (
    .PLUS(nd_aib39_ch5_x0y1),
    .MINUS(m1_ch5_aib[39])
   );

  aliasv xaliasv38_ch11 (
    .PLUS(nd_aib38_ch5_x0y1),
    .MINUS(m1_ch5_aib[38])
   );

  aliasv xaliasv37_ch11 (
    .PLUS(nd_aib37_ch5_x0y1),
    .MINUS(m1_ch5_aib[37])
   );

  aliasv xaliasv36_ch11 (
    .PLUS(nd_aib36_ch5_x0y1),
    .MINUS(m1_ch5_aib[36])
   );

  aliasv xaliasv35_ch11 (
    .PLUS(nd_aib35_ch5_x0y1),
    .MINUS(m1_ch5_aib[35])
   );

  aliasv xaliasv34_ch11 (
    .PLUS(nd_aib34_ch5_x0y1),
    .MINUS(m1_ch5_aib[34])
   );

  aliasv xaliasv33_ch11 (
    .PLUS(nd_aib33_ch5_x0y1),
    .MINUS(m1_ch5_aib[33])
   );

  aliasv xaliasv32_ch11 (
    .PLUS(nd_aib32_ch5_x0y1),
    .MINUS(m1_ch5_aib[32])
   );

  aliasv xaliasv31_ch11 (
    .PLUS(nd_aib31_ch5_x0y1),
    .MINUS(m1_ch5_aib[31])
   );

  aliasv xaliasv30_ch11 (
    .PLUS(nd_aib30_ch5_x0y1),
    .MINUS(m1_ch5_aib[30])
   );

  aliasv xaliasv29_ch11 (
    .PLUS(nd_aib29_ch5_x0y1),
    .MINUS(m1_ch5_aib[29])
   );

  aliasv xaliasv28_ch11 (
    .PLUS(nd_aib28_ch5_x0y1),
    .MINUS(m1_ch5_aib[28])
   );

  aliasv xaliasv27_ch11 (
    .PLUS(nd_aib27_ch5_x0y1),
    .MINUS(m1_ch5_aib[27])
   );

  aliasv xaliasv26_ch11 (
    .PLUS(nd_aib26_ch5_x0y1),
    .MINUS(m1_ch5_aib[26])
   );

  aliasv xaliasv25_ch11 (
    .PLUS(nd_aib25_ch5_x0y1),
    .MINUS(m1_ch5_aib[25])
   );

  aliasv xaliasv24_ch11 (
    .PLUS(nd_aib24_ch5_x0y1),
    .MINUS(m1_ch5_aib[24])
   );

  aliasv xaliasv23_ch11 (
    .PLUS(nd_aib23_ch5_x0y1),
    .MINUS(m1_ch5_aib[23])
   );

  aliasv xaliasv22_ch11 (
    .PLUS(nd_aib22_ch5_x0y1),
    .MINUS(m1_ch5_aib[22])
   );

  aliasv xaliasv21_ch11 (
    .PLUS(nd_aib21_ch5_x0y1),
    .MINUS(m1_ch5_aib[21])
   );

  aliasv xaliasv20_ch11 (
    .PLUS(nd_aib20_ch5_x0y1),
    .MINUS(m1_ch5_aib[20])
   );

  aliasv xaliasv19_ch11 (
    .PLUS(nd_aib19_ch5_x0y1),
    .MINUS(m1_ch5_aib[19])
   );

  aliasv xaliasv18_ch11 (
    .PLUS(nd_aib18_ch5_x0y1),
    .MINUS(m1_ch5_aib[18])
   );

  aliasv xaliasv17_ch11 (
    .PLUS(nd_aib17_ch5_x0y1),
    .MINUS(m1_ch5_aib[17])
   );

  aliasv xaliasv16_ch11 (
    .PLUS(nd_aib16_ch5_x0y1),
    .MINUS(m1_ch5_aib[16])
   );

  aliasv xaliasv15_ch11 (
    .PLUS(nd_aib15_ch5_x0y1),
    .MINUS(m1_ch5_aib[15])
   );

  aliasv xaliasv14_ch11 (
    .PLUS(nd_aib14_ch5_x0y1),
    .MINUS(m1_ch5_aib[14])
   );

  aliasv xaliasv13_ch11 (
    .PLUS(nd_aib13_ch5_x0y1),
    .MINUS(m1_ch5_aib[13])
   );

  aliasv xaliasv12_ch11 (
    .PLUS(nd_aib12_ch5_x0y1),
    .MINUS(m1_ch5_aib[12])
   );

  aliasv xaliasv11_ch11 (
    .PLUS(nd_aib11_ch5_x0y1),
    .MINUS(m1_ch5_aib[11])
   );

  aliasv xaliasv10_ch11 (
    .PLUS(nd_aib10_ch5_x0y1),
    .MINUS(m1_ch5_aib[10])
   );

  aliasv xaliasv9_ch11 (
    .PLUS(nd_aib9_ch5_x0y1),
    .MINUS(m1_ch5_aib[9])
   );

  aliasv xaliasv8_ch11 (
    .PLUS(nd_aib8_ch5_x0y1),
    .MINUS(m1_ch5_aib[8])
   );

  aliasv xaliasv7_ch11 (
    .PLUS(nd_aib7_ch5_x0y1),
    .MINUS(m1_ch5_aib[7])
   );

  aliasv xaliasv6_ch11 (
    .PLUS(nd_aib6_ch5_x0y1),
    .MINUS(m1_ch5_aib[6])
   );

  aliasv xaliasv5_ch11 (
    .PLUS(nd_aib5_ch5_x0y1),
    .MINUS(m1_ch5_aib[5])
   );

  aliasv xaliasv4_ch11 (
    .PLUS(nd_aib4_ch5_x0y1),
    .MINUS(m1_ch5_aib[4])
   );

  aliasv xaliasv3_ch11 (
    .PLUS(nd_aib3_ch5_x0y1),
    .MINUS(m1_ch5_aib[3])
   );

  aliasv xaliasv2_ch11 (
    .PLUS(nd_aib2_ch5_x0y1),
    .MINUS(m1_ch5_aib[2])
   );

  aliasv xaliasv1_ch11 (
    .PLUS(nd_aib1_ch5_x0y1),
    .MINUS(m1_ch5_aib[1])
   );

  aliasv xaliasv0_ch11 (
    .PLUS(nd_aib0_ch5_x0y1),
    .MINUS(m1_ch5_aib[0])
   );

// ## START OF ch12 ( ##
  aliasv xaliasv95_ch12 (
    .PLUS(nd_aib95_ch0_x0y2),
    .MINUS(m2_ch0_aib[95])
   );

  aliasv xaliasv94_ch12 (
    .PLUS(nd_aib94_ch0_x0y2),
    .MINUS(m2_ch0_aib[94])
   );

  aliasv xaliasv93_ch12 (
    .PLUS(nd_aib93_ch0_x0y2),
    .MINUS(m2_ch0_aib[93])
   );

  aliasv xaliasv92_ch12 (
    .PLUS(nd_aib92_ch0_x0y2),
    .MINUS(m2_ch0_aib[92])
   );

  aliasv xaliasv91_ch12 (
    .PLUS(nd_aib91_ch0_x0y2),
    .MINUS(m2_ch0_aib[91])
   );

  aliasv xaliasv90_ch12 (
    .PLUS(nd_aib90_ch0_x0y2),
    .MINUS(m2_ch0_aib[90])
   );

  aliasv xaliasv89_ch12 (
    .PLUS(nd_aib89_ch0_x0y2),
    .MINUS(m2_ch0_aib[89])
   );

  aliasv xaliasv88_ch12 (
    .PLUS(nd_aib88_ch0_x0y2),
    .MINUS(m2_ch0_aib[88])
   );

  aliasv xaliasv87_ch12 (
    .PLUS(nd_aib87_ch0_x0y2),
    .MINUS(m2_ch0_aib[87])
   );

  aliasv xaliasv86_ch12 (
    .PLUS(nd_aib86_ch0_x0y2),
    .MINUS(m2_ch0_aib[86])
   );

  aliasv xaliasv85_ch12 (
    .PLUS(nd_aib85_ch0_x0y2),
    .MINUS(m2_ch0_aib[85])
   );

  aliasv xaliasv84_ch12 (
    .PLUS(nd_aib84_ch0_x0y2),
    .MINUS(m2_ch0_aib[84])
   );

  aliasv xaliasv83_ch12 (
    .PLUS(nd_aib83_ch0_x0y2),
    .MINUS(m2_ch0_aib[83])
   );

  aliasv xaliasv82_ch12 (
    .PLUS(nd_aib82_ch0_x0y2),
    .MINUS(m2_ch0_aib[82])
   );

  aliasv xaliasv81_ch12 (
    .PLUS(nd_aib81_ch0_x0y2),
    .MINUS(m2_ch0_aib[81])
   );

  aliasv xaliasv80_ch12 (
    .PLUS(nd_aib80_ch0_x0y2),
    .MINUS(m2_ch0_aib[80])
   );

  aliasv xaliasv79_ch12 (
    .PLUS(nd_aib79_ch0_x0y2),
    .MINUS(m2_ch0_aib[79])
   );

  aliasv xaliasv78_ch12 (
    .PLUS(nd_aib78_ch0_x0y2),
    .MINUS(m2_ch0_aib[78])
   );

  aliasv xaliasv77_ch12 (
    .PLUS(nd_aib77_ch0_x0y2),
    .MINUS(m2_ch0_aib[77])
   );

  aliasv xaliasv76_ch12 (
    .PLUS(nd_aib76_ch0_x0y2),
    .MINUS(m2_ch0_aib[76])
   );

  aliasv xaliasv75_ch12 (
    .PLUS(nd_aib75_ch0_x0y2),
    .MINUS(m2_ch0_aib[75])
   );

  aliasv xaliasv74_ch12 (
    .PLUS(nd_aib74_ch0_x0y2),
    .MINUS(m2_ch0_aib[74])
   );

  aliasv xaliasv73_ch12 (
    .PLUS(nd_aib73_ch0_x0y2),
    .MINUS(m2_ch0_aib[73])
   );

  aliasv xaliasv72_ch12 (
    .PLUS(nd_aib72_ch0_x0y2),
    .MINUS(m2_ch0_aib[72])
   );

  aliasv xaliasv71_ch12 (
    .PLUS(nd_aib71_ch0_x0y2),
    .MINUS(m2_ch0_aib[71])
   );

  aliasv xaliasv70_ch12 (
    .PLUS(nd_aib70_ch0_x0y2),
    .MINUS(m2_ch0_aib[70])
   );

  aliasv xaliasv69_ch12 (
    .PLUS(nd_aib69_ch0_x0y2),
    .MINUS(m2_ch0_aib[69])
   );

  aliasv xaliasv68_ch12 (
    .PLUS(nd_aib68_ch0_x0y2),
    .MINUS(m2_ch0_aib[68])
   );

  aliasv xaliasv67_ch12 (
    .PLUS(nd_aib67_ch0_x0y2),
    .MINUS(m2_ch0_aib[67])
   );

  aliasv xaliasv66_ch12 (
    .PLUS(nd_aib66_ch0_x0y2),
    .MINUS(m2_ch0_aib[66])
   );

  aliasv xaliasv65_ch12 (
    .PLUS(nd_aib65_ch0_x0y2),
    .MINUS(m2_ch0_aib[65])
   );

  aliasv xaliasv64_ch12 (
    .PLUS(nd_aib64_ch0_x0y2),
    .MINUS(m2_ch0_aib[64])
   );

  aliasv xaliasv63_ch12 (
    .PLUS(nd_aib63_ch0_x0y2),
    .MINUS(m2_ch0_aib[63])
   );

  aliasv xaliasv62_ch12 (
    .PLUS(nd_aib62_ch0_x0y2),
    .MINUS(m2_ch0_aib[62])
   );

  aliasv xaliasv61_ch12 (
    .PLUS(nd_aib61_ch0_x0y2),
    .MINUS(m2_ch0_aib[61])
   );

  aliasv xaliasv60_ch12 (
    .PLUS(nd_aib60_ch0_x0y2),
    .MINUS(m2_ch0_aib[60])
   );

  aliasv xaliasv59_ch12 (
    .PLUS(nd_aib59_ch0_x0y2),
    .MINUS(m2_ch0_aib[59])
   );

  aliasv xaliasv58_ch12 (
    .PLUS(nd_aib58_ch0_x0y2),
    .MINUS(m2_ch0_aib[58])
   );

  aliasv xaliasv57_ch12 (
    .PLUS(nd_aib57_ch0_x0y2),
    .MINUS(m2_ch0_aib[57])
   );

  aliasv xaliasv56_ch12 (
    .PLUS(nd_aib56_ch0_x0y2),
    .MINUS(m2_ch0_aib[56])
   );

  aliasv xaliasv55_ch12 (
    .PLUS(nd_aib55_ch0_x0y2),
    .MINUS(m2_ch0_aib[55])
   );

  aliasv xaliasv54_ch12 (
    .PLUS(nd_aib54_ch0_x0y2),
    .MINUS(m2_ch0_aib[54])
   );

  aliasv xaliasv53_ch12 (
    .PLUS(nd_aib53_ch0_x0y2),
    .MINUS(m2_ch0_aib[53])
   );

  aliasv xaliasv52_ch12 (
    .PLUS(nd_aib52_ch0_x0y2),
    .MINUS(m2_ch0_aib[52])
   );

  aliasv xaliasv51_ch12 (
    .PLUS(nd_aib51_ch0_x0y2),
    .MINUS(m2_ch0_aib[51])
   );

  aliasv xaliasv50_ch12 (
    .PLUS(nd_aib50_ch0_x0y2),
    .MINUS(m2_ch0_aib[50])
   );

  aliasv xaliasv49_ch12 (
    .PLUS(nd_aib49_ch0_x0y2),
    .MINUS(m2_ch0_aib[49])
   );

  aliasv xaliasv48_ch12 (
    .PLUS(nd_aib48_ch0_x0y2),
    .MINUS(m2_ch0_aib[48])
   );

  aliasv xaliasv47_ch12 (
    .PLUS(nd_aib47_ch0_x0y2),
    .MINUS(m2_ch0_aib[47])
   );

  aliasv xaliasv46_ch12 (
    .PLUS(nd_aib46_ch0_x0y2),
    .MINUS(m2_ch0_aib[46])
   );

  aliasv xaliasv45_ch12 (
    .PLUS(nd_aib45_ch0_x0y2),
    .MINUS(m2_ch0_aib[45])
   );

  aliasv xaliasv44_ch12 (
    .PLUS(nd_aib44_ch0_x0y2),
    .MINUS(m2_ch0_aib[44])
   );

  aliasv xaliasv43_ch12 (
    .PLUS(nd_aib43_ch0_x0y2),
    .MINUS(m2_ch0_aib[43])
   );

  aliasv xaliasv42_ch12 (
    .PLUS(nd_aib42_ch0_x0y2),
    .MINUS(m2_ch0_aib[42])
   );

  aliasv xaliasv41_ch12 (
    .PLUS(nd_aib41_ch0_x0y2),
    .MINUS(m2_ch0_aib[41])
   );

  aliasv xaliasv40_ch12 (
    .PLUS(nd_aib40_ch0_x0y2),
    .MINUS(m2_ch0_aib[40])
   );

  aliasv xaliasv39_ch12 (
    .PLUS(nd_aib39_ch0_x0y2),
    .MINUS(m2_ch0_aib[39])
   );

  aliasv xaliasv38_ch12 (
    .PLUS(nd_aib38_ch0_x0y2),
    .MINUS(m2_ch0_aib[38])
   );

  aliasv xaliasv37_ch12 (
    .PLUS(nd_aib37_ch0_x0y2),
    .MINUS(m2_ch0_aib[37])
   );

  aliasv xaliasv36_ch12 (
    .PLUS(nd_aib36_ch0_x0y2),
    .MINUS(m2_ch0_aib[36])
   );

  aliasv xaliasv35_ch12 (
    .PLUS(nd_aib35_ch0_x0y2),
    .MINUS(m2_ch0_aib[35])
   );

  aliasv xaliasv34_ch12 (
    .PLUS(nd_aib34_ch0_x0y2),
    .MINUS(m2_ch0_aib[34])
   );

  aliasv xaliasv33_ch12 (
    .PLUS(nd_aib33_ch0_x0y2),
    .MINUS(m2_ch0_aib[33])
   );

  aliasv xaliasv32_ch12 (
    .PLUS(nd_aib32_ch0_x0y2),
    .MINUS(m2_ch0_aib[32])
   );

  aliasv xaliasv31_ch12 (
    .PLUS(nd_aib31_ch0_x0y2),
    .MINUS(m2_ch0_aib[31])
   );

  aliasv xaliasv30_ch12 (
    .PLUS(nd_aib30_ch0_x0y2),
    .MINUS(m2_ch0_aib[30])
   );

  aliasv xaliasv29_ch12 (
    .PLUS(nd_aib29_ch0_x0y2),
    .MINUS(m2_ch0_aib[29])
   );

  aliasv xaliasv28_ch12 (
    .PLUS(nd_aib28_ch0_x0y2),
    .MINUS(m2_ch0_aib[28])
   );

  aliasv xaliasv27_ch12 (
    .PLUS(nd_aib27_ch0_x0y2),
    .MINUS(m2_ch0_aib[27])
   );

  aliasv xaliasv26_ch12 (
    .PLUS(nd_aib26_ch0_x0y2),
    .MINUS(m2_ch0_aib[26])
   );

  aliasv xaliasv25_ch12 (
    .PLUS(nd_aib25_ch0_x0y2),
    .MINUS(m2_ch0_aib[25])
   );

  aliasv xaliasv24_ch12 (
    .PLUS(nd_aib24_ch0_x0y2),
    .MINUS(m2_ch0_aib[24])
   );

  aliasv xaliasv23_ch12 (
    .PLUS(nd_aib23_ch0_x0y2),
    .MINUS(m2_ch0_aib[23])
   );

  aliasv xaliasv22_ch12 (
    .PLUS(nd_aib22_ch0_x0y2),
    .MINUS(m2_ch0_aib[22])
   );

  aliasv xaliasv21_ch12 (
    .PLUS(nd_aib21_ch0_x0y2),
    .MINUS(m2_ch0_aib[21])
   );

  aliasv xaliasv20_ch12 (
    .PLUS(nd_aib20_ch0_x0y2),
    .MINUS(m2_ch0_aib[20])
   );

  aliasv xaliasv19_ch12 (
    .PLUS(nd_aib19_ch0_x0y2),
    .MINUS(m2_ch0_aib[19])
   );

  aliasv xaliasv18_ch12 (
    .PLUS(nd_aib18_ch0_x0y2),
    .MINUS(m2_ch0_aib[18])
   );

  aliasv xaliasv17_ch12 (
    .PLUS(nd_aib17_ch0_x0y2),
    .MINUS(m2_ch0_aib[17])
   );

  aliasv xaliasv16_ch12 (
    .PLUS(nd_aib16_ch0_x0y2),
    .MINUS(m2_ch0_aib[16])
   );

  aliasv xaliasv15_ch12 (
    .PLUS(nd_aib15_ch0_x0y2),
    .MINUS(m2_ch0_aib[15])
   );

  aliasv xaliasv14_ch12 (
    .PLUS(nd_aib14_ch0_x0y2),
    .MINUS(m2_ch0_aib[14])
   );

  aliasv xaliasv13_ch12 (
    .PLUS(nd_aib13_ch0_x0y2),
    .MINUS(m2_ch0_aib[13])
   );

  aliasv xaliasv12_ch12 (
    .PLUS(nd_aib12_ch0_x0y2),
    .MINUS(m2_ch0_aib[12])
   );

  aliasv xaliasv11_ch12 (
    .PLUS(nd_aib11_ch0_x0y2),
    .MINUS(m2_ch0_aib[11])
   );

  aliasv xaliasv10_ch12 (
    .PLUS(nd_aib10_ch0_x0y2),
    .MINUS(m2_ch0_aib[10])
   );

  aliasv xaliasv9_ch12 (
    .PLUS(nd_aib9_ch0_x0y2),
    .MINUS(m2_ch0_aib[9])
   );

  aliasv xaliasv8_ch12 (
    .PLUS(nd_aib8_ch0_x0y2),
    .MINUS(m2_ch0_aib[8])
   );

  aliasv xaliasv7_ch12 (
    .PLUS(nd_aib7_ch0_x0y2),
    .MINUS(m2_ch0_aib[7])
   );

  aliasv xaliasv6_ch12 (
    .PLUS(nd_aib6_ch0_x0y2),
    .MINUS(m2_ch0_aib[6])
   );

  aliasv xaliasv5_ch12 (
    .PLUS(nd_aib5_ch0_x0y2),
    .MINUS(m2_ch0_aib[5])
   );

  aliasv xaliasv4_ch12 (
    .PLUS(nd_aib4_ch0_x0y2),
    .MINUS(m2_ch0_aib[4])
   );

  aliasv xaliasv3_ch12 (
    .PLUS(nd_aib3_ch0_x0y2),
    .MINUS(m2_ch0_aib[3])
   );

  aliasv xaliasv2_ch12 (
    .PLUS(nd_aib2_ch0_x0y2),
    .MINUS(m2_ch0_aib[2])
   );

  aliasv xaliasv1_ch12 (
    .PLUS(nd_aib1_ch0_x0y2),
    .MINUS(m2_ch0_aib[1])
   );

  aliasv xaliasv0_ch12 (
    .PLUS(nd_aib0_ch0_x0y2),
    .MINUS(m2_ch0_aib[0])
   );

// ## START OF ch13 ( ##
  aliasv xaliasv95_ch13 (
    .PLUS(nd_aib95_ch1_x0y2),
    .MINUS(m2_ch1_aib[95])
   );

  aliasv xaliasv94_ch13 (
    .PLUS(nd_aib94_ch1_x0y2),
    .MINUS(m2_ch1_aib[94])
   );

  aliasv xaliasv93_ch13 (
    .PLUS(nd_aib93_ch1_x0y2),
    .MINUS(m2_ch1_aib[93])
   );

  aliasv xaliasv92_ch13 (
    .PLUS(nd_aib92_ch1_x0y2),
    .MINUS(m2_ch1_aib[92])
   );

  aliasv xaliasv91_ch13 (
    .PLUS(nd_aib91_ch1_x0y2),
    .MINUS(m2_ch1_aib[91])
   );

  aliasv xaliasv90_ch13 (
    .PLUS(nd_aib90_ch1_x0y2),
    .MINUS(m2_ch1_aib[90])
   );

  aliasv xaliasv89_ch13 (
    .PLUS(nd_aib89_ch1_x0y2),
    .MINUS(m2_ch1_aib[89])
   );

  aliasv xaliasv88_ch13 (
    .PLUS(nd_aib88_ch1_x0y2),
    .MINUS(m2_ch1_aib[88])
   );

  aliasv xaliasv87_ch13 (
    .PLUS(nd_aib87_ch1_x0y2),
    .MINUS(m2_ch1_aib[87])
   );

  aliasv xaliasv86_ch13 (
    .PLUS(nd_aib86_ch1_x0y2),
    .MINUS(m2_ch1_aib[86])
   );

  aliasv xaliasv85_ch13 (
    .PLUS(nd_aib85_ch1_x0y2),
    .MINUS(m2_ch1_aib[85])
   );

  aliasv xaliasv84_ch13 (
    .PLUS(nd_aib84_ch1_x0y2),
    .MINUS(m2_ch1_aib[84])
   );

  aliasv xaliasv83_ch13 (
    .PLUS(nd_aib83_ch1_x0y2),
    .MINUS(m2_ch1_aib[83])
   );

  aliasv xaliasv82_ch13 (
    .PLUS(nd_aib82_ch1_x0y2),
    .MINUS(m2_ch1_aib[82])
   );

  aliasv xaliasv81_ch13 (
    .PLUS(nd_aib81_ch1_x0y2),
    .MINUS(m2_ch1_aib[81])
   );

  aliasv xaliasv80_ch13 (
    .PLUS(nd_aib80_ch1_x0y2),
    .MINUS(m2_ch1_aib[80])
   );

  aliasv xaliasv79_ch13 (
    .PLUS(nd_aib79_ch1_x0y2),
    .MINUS(m2_ch1_aib[79])
   );

  aliasv xaliasv78_ch13 (
    .PLUS(nd_aib78_ch1_x0y2),
    .MINUS(m2_ch1_aib[78])
   );

  aliasv xaliasv77_ch13 (
    .PLUS(nd_aib77_ch1_x0y2),
    .MINUS(m2_ch1_aib[77])
   );

  aliasv xaliasv76_ch13 (
    .PLUS(nd_aib76_ch1_x0y2),
    .MINUS(m2_ch1_aib[76])
   );

  aliasv xaliasv75_ch13 (
    .PLUS(nd_aib75_ch1_x0y2),
    .MINUS(m2_ch1_aib[75])
   );

  aliasv xaliasv74_ch13 (
    .PLUS(nd_aib74_ch1_x0y2),
    .MINUS(m2_ch1_aib[74])
   );

  aliasv xaliasv73_ch13 (
    .PLUS(nd_aib73_ch1_x0y2),
    .MINUS(m2_ch1_aib[73])
   );

  aliasv xaliasv72_ch13 (
    .PLUS(nd_aib72_ch1_x0y2),
    .MINUS(m2_ch1_aib[72])
   );

  aliasv xaliasv71_ch13 (
    .PLUS(nd_aib71_ch1_x0y2),
    .MINUS(m2_ch1_aib[71])
   );

  aliasv xaliasv70_ch13 (
    .PLUS(nd_aib70_ch1_x0y2),
    .MINUS(m2_ch1_aib[70])
   );

  aliasv xaliasv69_ch13 (
    .PLUS(nd_aib69_ch1_x0y2),
    .MINUS(m2_ch1_aib[69])
   );

  aliasv xaliasv68_ch13 (
    .PLUS(nd_aib68_ch1_x0y2),
    .MINUS(m2_ch1_aib[68])
   );

  aliasv xaliasv67_ch13 (
    .PLUS(nd_aib67_ch1_x0y2),
    .MINUS(m2_ch1_aib[67])
   );

  aliasv xaliasv66_ch13 (
    .PLUS(nd_aib66_ch1_x0y2),
    .MINUS(m2_ch1_aib[66])
   );

  aliasv xaliasv65_ch13 (
    .PLUS(nd_aib65_ch1_x0y2),
    .MINUS(m2_ch1_aib[65])
   );

  aliasv xaliasv64_ch13 (
    .PLUS(nd_aib64_ch1_x0y2),
    .MINUS(m2_ch1_aib[64])
   );

  aliasv xaliasv63_ch13 (
    .PLUS(nd_aib63_ch1_x0y2),
    .MINUS(m2_ch1_aib[63])
   );

  aliasv xaliasv62_ch13 (
    .PLUS(nd_aib62_ch1_x0y2),
    .MINUS(m2_ch1_aib[62])
   );

  aliasv xaliasv61_ch13 (
    .PLUS(nd_aib61_ch1_x0y2),
    .MINUS(m2_ch1_aib[61])
   );

  aliasv xaliasv60_ch13 (
    .PLUS(nd_aib60_ch1_x0y2),
    .MINUS(m2_ch1_aib[60])
   );

  aliasv xaliasv59_ch13 (
    .PLUS(nd_aib59_ch1_x0y2),
    .MINUS(m2_ch1_aib[59])
   );

  aliasv xaliasv58_ch13 (
    .PLUS(nd_aib58_ch1_x0y2),
    .MINUS(m2_ch1_aib[58])
   );

  aliasv xaliasv57_ch13 (
    .PLUS(nd_aib57_ch1_x0y2),
    .MINUS(m2_ch1_aib[57])
   );

  aliasv xaliasv56_ch13 (
    .PLUS(nd_aib56_ch1_x0y2),
    .MINUS(m2_ch1_aib[56])
   );

  aliasv xaliasv55_ch13 (
    .PLUS(nd_aib55_ch1_x0y2),
    .MINUS(m2_ch1_aib[55])
   );

  aliasv xaliasv54_ch13 (
    .PLUS(nd_aib54_ch1_x0y2),
    .MINUS(m2_ch1_aib[54])
   );

  aliasv xaliasv53_ch13 (
    .PLUS(nd_aib53_ch1_x0y2),
    .MINUS(m2_ch1_aib[53])
   );

  aliasv xaliasv52_ch13 (
    .PLUS(nd_aib52_ch1_x0y2),
    .MINUS(m2_ch1_aib[52])
   );

  aliasv xaliasv51_ch13 (
    .PLUS(nd_aib51_ch1_x0y2),
    .MINUS(m2_ch1_aib[51])
   );

  aliasv xaliasv50_ch13 (
    .PLUS(nd_aib50_ch1_x0y2),
    .MINUS(m2_ch1_aib[50])
   );

  aliasv xaliasv49_ch13 (
    .PLUS(nd_aib49_ch1_x0y2),
    .MINUS(m2_ch1_aib[49])
   );

  aliasv xaliasv48_ch13 (
    .PLUS(nd_aib48_ch1_x0y2),
    .MINUS(m2_ch1_aib[48])
   );

  aliasv xaliasv47_ch13 (
    .PLUS(nd_aib47_ch1_x0y2),
    .MINUS(m2_ch1_aib[47])
   );

  aliasv xaliasv46_ch13 (
    .PLUS(nd_aib46_ch1_x0y2),
    .MINUS(m2_ch1_aib[46])
   );

  aliasv xaliasv45_ch13 (
    .PLUS(nd_aib45_ch1_x0y2),
    .MINUS(m2_ch1_aib[45])
   );

  aliasv xaliasv44_ch13 (
    .PLUS(nd_aib44_ch1_x0y2),
    .MINUS(m2_ch1_aib[44])
   );

  aliasv xaliasv43_ch13 (
    .PLUS(nd_aib43_ch1_x0y2),
    .MINUS(m2_ch1_aib[43])
   );

  aliasv xaliasv42_ch13 (
    .PLUS(nd_aib42_ch1_x0y2),
    .MINUS(m2_ch1_aib[42])
   );

  aliasv xaliasv41_ch13 (
    .PLUS(nd_aib41_ch1_x0y2),
    .MINUS(m2_ch1_aib[41])
   );

  aliasv xaliasv40_ch13 (
    .PLUS(nd_aib40_ch1_x0y2),
    .MINUS(m2_ch1_aib[40])
   );

  aliasv xaliasv39_ch13 (
    .PLUS(nd_aib39_ch1_x0y2),
    .MINUS(m2_ch1_aib[39])
   );

  aliasv xaliasv38_ch13 (
    .PLUS(nd_aib38_ch1_x0y2),
    .MINUS(m2_ch1_aib[38])
   );

  aliasv xaliasv37_ch13 (
    .PLUS(nd_aib37_ch1_x0y2),
    .MINUS(m2_ch1_aib[37])
   );

  aliasv xaliasv36_ch13 (
    .PLUS(nd_aib36_ch1_x0y2),
    .MINUS(m2_ch1_aib[36])
   );

  aliasv xaliasv35_ch13 (
    .PLUS(nd_aib35_ch1_x0y2),
    .MINUS(m2_ch1_aib[35])
   );

  aliasv xaliasv34_ch13 (
    .PLUS(nd_aib34_ch1_x0y2),
    .MINUS(m2_ch1_aib[34])
   );

  aliasv xaliasv33_ch13 (
    .PLUS(nd_aib33_ch1_x0y2),
    .MINUS(m2_ch1_aib[33])
   );

  aliasv xaliasv32_ch13 (
    .PLUS(nd_aib32_ch1_x0y2),
    .MINUS(m2_ch1_aib[32])
   );

  aliasv xaliasv31_ch13 (
    .PLUS(nd_aib31_ch1_x0y2),
    .MINUS(m2_ch1_aib[31])
   );

  aliasv xaliasv30_ch13 (
    .PLUS(nd_aib30_ch1_x0y2),
    .MINUS(m2_ch1_aib[30])
   );

  aliasv xaliasv29_ch13 (
    .PLUS(nd_aib29_ch1_x0y2),
    .MINUS(m2_ch1_aib[29])
   );

  aliasv xaliasv28_ch13 (
    .PLUS(nd_aib28_ch1_x0y2),
    .MINUS(m2_ch1_aib[28])
   );

  aliasv xaliasv27_ch13 (
    .PLUS(nd_aib27_ch1_x0y2),
    .MINUS(m2_ch1_aib[27])
   );

  aliasv xaliasv26_ch13 (
    .PLUS(nd_aib26_ch1_x0y2),
    .MINUS(m2_ch1_aib[26])
   );

  aliasv xaliasv25_ch13 (
    .PLUS(nd_aib25_ch1_x0y2),
    .MINUS(m2_ch1_aib[25])
   );

  aliasv xaliasv24_ch13 (
    .PLUS(nd_aib24_ch1_x0y2),
    .MINUS(m2_ch1_aib[24])
   );

  aliasv xaliasv23_ch13 (
    .PLUS(nd_aib23_ch1_x0y2),
    .MINUS(m2_ch1_aib[23])
   );

  aliasv xaliasv22_ch13 (
    .PLUS(nd_aib22_ch1_x0y2),
    .MINUS(m2_ch1_aib[22])
   );

  aliasv xaliasv21_ch13 (
    .PLUS(nd_aib21_ch1_x0y2),
    .MINUS(m2_ch1_aib[21])
   );

  aliasv xaliasv20_ch13 (
    .PLUS(nd_aib20_ch1_x0y2),
    .MINUS(m2_ch1_aib[20])
   );

  aliasv xaliasv19_ch13 (
    .PLUS(nd_aib19_ch1_x0y2),
    .MINUS(m2_ch1_aib[19])
   );

  aliasv xaliasv18_ch13 (
    .PLUS(nd_aib18_ch1_x0y2),
    .MINUS(m2_ch1_aib[18])
   );

  aliasv xaliasv17_ch13 (
    .PLUS(nd_aib17_ch1_x0y2),
    .MINUS(m2_ch1_aib[17])
   );

  aliasv xaliasv16_ch13 (
    .PLUS(nd_aib16_ch1_x0y2),
    .MINUS(m2_ch1_aib[16])
   );

  aliasv xaliasv15_ch13 (
    .PLUS(nd_aib15_ch1_x0y2),
    .MINUS(m2_ch1_aib[15])
   );

  aliasv xaliasv14_ch13 (
    .PLUS(nd_aib14_ch1_x0y2),
    .MINUS(m2_ch1_aib[14])
   );

  aliasv xaliasv13_ch13 (
    .PLUS(nd_aib13_ch1_x0y2),
    .MINUS(m2_ch1_aib[13])
   );

  aliasv xaliasv12_ch13 (
    .PLUS(nd_aib12_ch1_x0y2),
    .MINUS(m2_ch1_aib[12])
   );

  aliasv xaliasv11_ch13 (
    .PLUS(nd_aib11_ch1_x0y2),
    .MINUS(m2_ch1_aib[11])
   );

  aliasv xaliasv10_ch13 (
    .PLUS(nd_aib10_ch1_x0y2),
    .MINUS(m2_ch1_aib[10])
   );

  aliasv xaliasv9_ch13 (
    .PLUS(nd_aib9_ch1_x0y2),
    .MINUS(m2_ch1_aib[9])
   );

  aliasv xaliasv8_ch13 (
    .PLUS(nd_aib8_ch1_x0y2),
    .MINUS(m2_ch1_aib[8])
   );

  aliasv xaliasv7_ch13 (
    .PLUS(nd_aib7_ch1_x0y2),
    .MINUS(m2_ch1_aib[7])
   );

  aliasv xaliasv6_ch13 (
    .PLUS(nd_aib6_ch1_x0y2),
    .MINUS(m2_ch1_aib[6])
   );

  aliasv xaliasv5_ch13 (
    .PLUS(nd_aib5_ch1_x0y2),
    .MINUS(m2_ch1_aib[5])
   );

  aliasv xaliasv4_ch13 (
    .PLUS(nd_aib4_ch1_x0y2),
    .MINUS(m2_ch1_aib[4])
   );

  aliasv xaliasv3_ch13 (
    .PLUS(nd_aib3_ch1_x0y2),
    .MINUS(m2_ch1_aib[3])
   );

  aliasv xaliasv2_ch13 (
    .PLUS(nd_aib2_ch1_x0y2),
    .MINUS(m2_ch1_aib[2])
   );

  aliasv xaliasv1_ch13 (
    .PLUS(nd_aib1_ch1_x0y2),
    .MINUS(m2_ch1_aib[1])
   );

  aliasv xaliasv0_ch13 (
    .PLUS(nd_aib0_ch1_x0y2),
    .MINUS(m2_ch1_aib[0])
   );

// ## START OF ch14 ( ##
  aliasv xaliasv95_ch14 (
    .PLUS(nd_aib95_ch2_x0y2),
    .MINUS(m2_ch2_aib[95])
   );

  aliasv xaliasv94_ch14 (
    .PLUS(nd_aib94_ch2_x0y2),
    .MINUS(m2_ch2_aib[94])
   );

  aliasv xaliasv93_ch14 (
    .PLUS(nd_aib93_ch2_x0y2),
    .MINUS(m2_ch2_aib[93])
   );

  aliasv xaliasv92_ch14 (
    .PLUS(nd_aib92_ch2_x0y2),
    .MINUS(m2_ch2_aib[92])
   );

  aliasv xaliasv91_ch14 (
    .PLUS(nd_aib91_ch2_x0y2),
    .MINUS(m2_ch2_aib[91])
   );

  aliasv xaliasv90_ch14 (
    .PLUS(nd_aib90_ch2_x0y2),
    .MINUS(m2_ch2_aib[90])
   );

  aliasv xaliasv89_ch14 (
    .PLUS(nd_aib89_ch2_x0y2),
    .MINUS(m2_ch2_aib[89])
   );

  aliasv xaliasv88_ch14 (
    .PLUS(nd_aib88_ch2_x0y2),
    .MINUS(m2_ch2_aib[88])
   );

  aliasv xaliasv87_ch14 (
    .PLUS(nd_aib87_ch2_x0y2),
    .MINUS(m2_ch2_aib[87])
   );

  aliasv xaliasv86_ch14 (
    .PLUS(nd_aib86_ch2_x0y2),
    .MINUS(m2_ch2_aib[86])
   );

  aliasv xaliasv85_ch14 (
    .PLUS(nd_aib85_ch2_x0y2),
    .MINUS(m2_ch2_aib[85])
   );

  aliasv xaliasv84_ch14 (
    .PLUS(nd_aib84_ch2_x0y2),
    .MINUS(m2_ch2_aib[84])
   );

  aliasv xaliasv83_ch14 (
    .PLUS(nd_aib83_ch2_x0y2),
    .MINUS(m2_ch2_aib[83])
   );

  aliasv xaliasv82_ch14 (
    .PLUS(nd_aib82_ch2_x0y2),
    .MINUS(m2_ch2_aib[82])
   );

  aliasv xaliasv81_ch14 (
    .PLUS(nd_aib81_ch2_x0y2),
    .MINUS(m2_ch2_aib[81])
   );

  aliasv xaliasv80_ch14 (
    .PLUS(nd_aib80_ch2_x0y2),
    .MINUS(m2_ch2_aib[80])
   );

  aliasv xaliasv79_ch14 (
    .PLUS(nd_aib79_ch2_x0y2),
    .MINUS(m2_ch2_aib[79])
   );

  aliasv xaliasv78_ch14 (
    .PLUS(nd_aib78_ch2_x0y2),
    .MINUS(m2_ch2_aib[78])
   );

  aliasv xaliasv77_ch14 (
    .PLUS(nd_aib77_ch2_x0y2),
    .MINUS(m2_ch2_aib[77])
   );

  aliasv xaliasv76_ch14 (
    .PLUS(nd_aib76_ch2_x0y2),
    .MINUS(m2_ch2_aib[76])
   );

  aliasv xaliasv75_ch14 (
    .PLUS(nd_aib75_ch2_x0y2),
    .MINUS(m2_ch2_aib[75])
   );

  aliasv xaliasv74_ch14 (
    .PLUS(nd_aib74_ch2_x0y2),
    .MINUS(m2_ch2_aib[74])
   );

  aliasv xaliasv73_ch14 (
    .PLUS(nd_aib73_ch2_x0y2),
    .MINUS(m2_ch2_aib[73])
   );

  aliasv xaliasv72_ch14 (
    .PLUS(nd_aib72_ch2_x0y2),
    .MINUS(m2_ch2_aib[72])
   );

  aliasv xaliasv71_ch14 (
    .PLUS(nd_aib71_ch2_x0y2),
    .MINUS(m2_ch2_aib[71])
   );

  aliasv xaliasv70_ch14 (
    .PLUS(nd_aib70_ch2_x0y2),
    .MINUS(m2_ch2_aib[70])
   );

  aliasv xaliasv69_ch14 (
    .PLUS(nd_aib69_ch2_x0y2),
    .MINUS(m2_ch2_aib[69])
   );

  aliasv xaliasv68_ch14 (
    .PLUS(nd_aib68_ch2_x0y2),
    .MINUS(m2_ch2_aib[68])
   );

  aliasv xaliasv67_ch14 (
    .PLUS(nd_aib67_ch2_x0y2),
    .MINUS(m2_ch2_aib[67])
   );

  aliasv xaliasv66_ch14 (
    .PLUS(nd_aib66_ch2_x0y2),
    .MINUS(m2_ch2_aib[66])
   );

  aliasv xaliasv65_ch14 (
    .PLUS(nd_aib65_ch2_x0y2),
    .MINUS(m2_ch2_aib[65])
   );

  aliasv xaliasv64_ch14 (
    .PLUS(nd_aib64_ch2_x0y2),
    .MINUS(m2_ch2_aib[64])
   );

  aliasv xaliasv63_ch14 (
    .PLUS(nd_aib63_ch2_x0y2),
    .MINUS(m2_ch2_aib[63])
   );

  aliasv xaliasv62_ch14 (
    .PLUS(nd_aib62_ch2_x0y2),
    .MINUS(m2_ch2_aib[62])
   );

  aliasv xaliasv61_ch14 (
    .PLUS(nd_aib61_ch2_x0y2),
    .MINUS(m2_ch2_aib[61])
   );

  aliasv xaliasv60_ch14 (
    .PLUS(nd_aib60_ch2_x0y2),
    .MINUS(m2_ch2_aib[60])
   );

  aliasv xaliasv59_ch14 (
    .PLUS(nd_aib59_ch2_x0y2),
    .MINUS(m2_ch2_aib[59])
   );

  aliasv xaliasv58_ch14 (
    .PLUS(nd_aib58_ch2_x0y2),
    .MINUS(m2_ch2_aib[58])
   );

  aliasv xaliasv57_ch14 (
    .PLUS(nd_aib57_ch2_x0y2),
    .MINUS(m2_ch2_aib[57])
   );

  aliasv xaliasv56_ch14 (
    .PLUS(nd_aib56_ch2_x0y2),
    .MINUS(m2_ch2_aib[56])
   );

  aliasv xaliasv55_ch14 (
    .PLUS(nd_aib55_ch2_x0y2),
    .MINUS(m2_ch2_aib[55])
   );

  aliasv xaliasv54_ch14 (
    .PLUS(nd_aib54_ch2_x0y2),
    .MINUS(m2_ch2_aib[54])
   );

  aliasv xaliasv53_ch14 (
    .PLUS(nd_aib53_ch2_x0y2),
    .MINUS(m2_ch2_aib[53])
   );

  aliasv xaliasv52_ch14 (
    .PLUS(nd_aib52_ch2_x0y2),
    .MINUS(m2_ch2_aib[52])
   );

  aliasv xaliasv51_ch14 (
    .PLUS(nd_aib51_ch2_x0y2),
    .MINUS(m2_ch2_aib[51])
   );

  aliasv xaliasv50_ch14 (
    .PLUS(nd_aib50_ch2_x0y2),
    .MINUS(m2_ch2_aib[50])
   );

  aliasv xaliasv49_ch14 (
    .PLUS(nd_aib49_ch2_x0y2),
    .MINUS(m2_ch2_aib[49])
   );

  aliasv xaliasv48_ch14 (
    .PLUS(nd_aib48_ch2_x0y2),
    .MINUS(m2_ch2_aib[48])
   );

  aliasv xaliasv47_ch14 (
    .PLUS(nd_aib47_ch2_x0y2),
    .MINUS(m2_ch2_aib[47])
   );

  aliasv xaliasv46_ch14 (
    .PLUS(nd_aib46_ch2_x0y2),
    .MINUS(m2_ch2_aib[46])
   );

  aliasv xaliasv45_ch14 (
    .PLUS(nd_aib45_ch2_x0y2),
    .MINUS(m2_ch2_aib[45])
   );

  aliasv xaliasv44_ch14 (
    .PLUS(nd_aib44_ch2_x0y2),
    .MINUS(m2_ch2_aib[44])
   );

  aliasv xaliasv43_ch14 (
    .PLUS(nd_aib43_ch2_x0y2),
    .MINUS(m2_ch2_aib[43])
   );

  aliasv xaliasv42_ch14 (
    .PLUS(nd_aib42_ch2_x0y2),
    .MINUS(m2_ch2_aib[42])
   );

  aliasv xaliasv41_ch14 (
    .PLUS(nd_aib41_ch2_x0y2),
    .MINUS(m2_ch2_aib[41])
   );

  aliasv xaliasv40_ch14 (
    .PLUS(nd_aib40_ch2_x0y2),
    .MINUS(m2_ch2_aib[40])
   );

  aliasv xaliasv39_ch14 (
    .PLUS(nd_aib39_ch2_x0y2),
    .MINUS(m2_ch2_aib[39])
   );

  aliasv xaliasv38_ch14 (
    .PLUS(nd_aib38_ch2_x0y2),
    .MINUS(m2_ch2_aib[38])
   );

  aliasv xaliasv37_ch14 (
    .PLUS(nd_aib37_ch2_x0y2),
    .MINUS(m2_ch2_aib[37])
   );

  aliasv xaliasv36_ch14 (
    .PLUS(nd_aib36_ch2_x0y2),
    .MINUS(m2_ch2_aib[36])
   );

  aliasv xaliasv35_ch14 (
    .PLUS(nd_aib35_ch2_x0y2),
    .MINUS(m2_ch2_aib[35])
   );

  aliasv xaliasv34_ch14 (
    .PLUS(nd_aib34_ch2_x0y2),
    .MINUS(m2_ch2_aib[34])
   );

  aliasv xaliasv33_ch14 (
    .PLUS(nd_aib33_ch2_x0y2),
    .MINUS(m2_ch2_aib[33])
   );

  aliasv xaliasv32_ch14 (
    .PLUS(nd_aib32_ch2_x0y2),
    .MINUS(m2_ch2_aib[32])
   );

  aliasv xaliasv31_ch14 (
    .PLUS(nd_aib31_ch2_x0y2),
    .MINUS(m2_ch2_aib[31])
   );

  aliasv xaliasv30_ch14 (
    .PLUS(nd_aib30_ch2_x0y2),
    .MINUS(m2_ch2_aib[30])
   );

  aliasv xaliasv29_ch14 (
    .PLUS(nd_aib29_ch2_x0y2),
    .MINUS(m2_ch2_aib[29])
   );

  aliasv xaliasv28_ch14 (
    .PLUS(nd_aib28_ch2_x0y2),
    .MINUS(m2_ch2_aib[28])
   );

  aliasv xaliasv27_ch14 (
    .PLUS(nd_aib27_ch2_x0y2),
    .MINUS(m2_ch2_aib[27])
   );

  aliasv xaliasv26_ch14 (
    .PLUS(nd_aib26_ch2_x0y2),
    .MINUS(m2_ch2_aib[26])
   );

  aliasv xaliasv25_ch14 (
    .PLUS(nd_aib25_ch2_x0y2),
    .MINUS(m2_ch2_aib[25])
   );

  aliasv xaliasv24_ch14 (
    .PLUS(nd_aib24_ch2_x0y2),
    .MINUS(m2_ch2_aib[24])
   );

  aliasv xaliasv23_ch14 (
    .PLUS(nd_aib23_ch2_x0y2),
    .MINUS(m2_ch2_aib[23])
   );

  aliasv xaliasv22_ch14 (
    .PLUS(nd_aib22_ch2_x0y2),
    .MINUS(m2_ch2_aib[22])
   );

  aliasv xaliasv21_ch14 (
    .PLUS(nd_aib21_ch2_x0y2),
    .MINUS(m2_ch2_aib[21])
   );

  aliasv xaliasv20_ch14 (
    .PLUS(nd_aib20_ch2_x0y2),
    .MINUS(m2_ch2_aib[20])
   );

  aliasv xaliasv19_ch14 (
    .PLUS(nd_aib19_ch2_x0y2),
    .MINUS(m2_ch2_aib[19])
   );

  aliasv xaliasv18_ch14 (
    .PLUS(nd_aib18_ch2_x0y2),
    .MINUS(m2_ch2_aib[18])
   );

  aliasv xaliasv17_ch14 (
    .PLUS(nd_aib17_ch2_x0y2),
    .MINUS(m2_ch2_aib[17])
   );

  aliasv xaliasv16_ch14 (
    .PLUS(nd_aib16_ch2_x0y2),
    .MINUS(m2_ch2_aib[16])
   );

  aliasv xaliasv15_ch14 (
    .PLUS(nd_aib15_ch2_x0y2),
    .MINUS(m2_ch2_aib[15])
   );

  aliasv xaliasv14_ch14 (
    .PLUS(nd_aib14_ch2_x0y2),
    .MINUS(m2_ch2_aib[14])
   );

  aliasv xaliasv13_ch14 (
    .PLUS(nd_aib13_ch2_x0y2),
    .MINUS(m2_ch2_aib[13])
   );

  aliasv xaliasv12_ch14 (
    .PLUS(nd_aib12_ch2_x0y2),
    .MINUS(m2_ch2_aib[12])
   );

  aliasv xaliasv11_ch14 (
    .PLUS(nd_aib11_ch2_x0y2),
    .MINUS(m2_ch2_aib[11])
   );

  aliasv xaliasv10_ch14 (
    .PLUS(nd_aib10_ch2_x0y2),
    .MINUS(m2_ch2_aib[10])
   );

  aliasv xaliasv9_ch14 (
    .PLUS(nd_aib9_ch2_x0y2),
    .MINUS(m2_ch2_aib[9])
   );

  aliasv xaliasv8_ch14 (
    .PLUS(nd_aib8_ch2_x0y2),
    .MINUS(m2_ch2_aib[8])
   );

  aliasv xaliasv7_ch14 (
    .PLUS(nd_aib7_ch2_x0y2),
    .MINUS(m2_ch2_aib[7])
   );

  aliasv xaliasv6_ch14 (
    .PLUS(nd_aib6_ch2_x0y2),
    .MINUS(m2_ch2_aib[6])
   );

  aliasv xaliasv5_ch14 (
    .PLUS(nd_aib5_ch2_x0y2),
    .MINUS(m2_ch2_aib[5])
   );

  aliasv xaliasv4_ch14 (
    .PLUS(nd_aib4_ch2_x0y2),
    .MINUS(m2_ch2_aib[4])
   );

  aliasv xaliasv3_ch14 (
    .PLUS(nd_aib3_ch2_x0y2),
    .MINUS(m2_ch2_aib[3])
   );

  aliasv xaliasv2_ch14 (
    .PLUS(nd_aib2_ch2_x0y2),
    .MINUS(m2_ch2_aib[2])
   );

  aliasv xaliasv1_ch14 (
    .PLUS(nd_aib1_ch2_x0y2),
    .MINUS(m2_ch2_aib[1])
   );

  aliasv xaliasv0_ch14 (
    .PLUS(nd_aib0_ch2_x0y2),
    .MINUS(m2_ch2_aib[0])
   );

// ## START OF ch15 ( ##
  aliasv xaliasv95_ch15 (
    .PLUS(nd_aib95_ch3_x0y2),
    .MINUS(m2_ch3_aib[95])
   );

  aliasv xaliasv94_ch15 (
    .PLUS(nd_aib94_ch3_x0y2),
    .MINUS(m2_ch3_aib[94])
   );

  aliasv xaliasv93_ch15 (
    .PLUS(nd_aib93_ch3_x0y2),
    .MINUS(m2_ch3_aib[93])
   );

  aliasv xaliasv92_ch15 (
    .PLUS(nd_aib92_ch3_x0y2),
    .MINUS(m2_ch3_aib[92])
   );

  aliasv xaliasv91_ch15 (
    .PLUS(nd_aib91_ch3_x0y2),
    .MINUS(m2_ch3_aib[91])
   );

  aliasv xaliasv90_ch15 (
    .PLUS(nd_aib90_ch3_x0y2),
    .MINUS(m2_ch3_aib[90])
   );

  aliasv xaliasv89_ch15 (
    .PLUS(nd_aib89_ch3_x0y2),
    .MINUS(m2_ch3_aib[89])
   );

  aliasv xaliasv88_ch15 (
    .PLUS(nd_aib88_ch3_x0y2),
    .MINUS(m2_ch3_aib[88])
   );

  aliasv xaliasv87_ch15 (
    .PLUS(nd_aib87_ch3_x0y2),
    .MINUS(m2_ch3_aib[87])
   );

  aliasv xaliasv86_ch15 (
    .PLUS(nd_aib86_ch3_x0y2),
    .MINUS(m2_ch3_aib[86])
   );

  aliasv xaliasv85_ch15 (
    .PLUS(nd_aib85_ch3_x0y2),
    .MINUS(m2_ch3_aib[85])
   );

  aliasv xaliasv84_ch15 (
    .PLUS(nd_aib84_ch3_x0y2),
    .MINUS(m2_ch3_aib[84])
   );

  aliasv xaliasv83_ch15 (
    .PLUS(nd_aib83_ch3_x0y2),
    .MINUS(m2_ch3_aib[83])
   );

  aliasv xaliasv82_ch15 (
    .PLUS(nd_aib82_ch3_x0y2),
    .MINUS(m2_ch3_aib[82])
   );

  aliasv xaliasv81_ch15 (
    .PLUS(nd_aib81_ch3_x0y2),
    .MINUS(m2_ch3_aib[81])
   );

  aliasv xaliasv80_ch15 (
    .PLUS(nd_aib80_ch3_x0y2),
    .MINUS(m2_ch3_aib[80])
   );

  aliasv xaliasv79_ch15 (
    .PLUS(nd_aib79_ch3_x0y2),
    .MINUS(m2_ch3_aib[79])
   );

  aliasv xaliasv78_ch15 (
    .PLUS(nd_aib78_ch3_x0y2),
    .MINUS(m2_ch3_aib[78])
   );

  aliasv xaliasv77_ch15 (
    .PLUS(nd_aib77_ch3_x0y2),
    .MINUS(m2_ch3_aib[77])
   );

  aliasv xaliasv76_ch15 (
    .PLUS(nd_aib76_ch3_x0y2),
    .MINUS(m2_ch3_aib[76])
   );

  aliasv xaliasv75_ch15 (
    .PLUS(nd_aib75_ch3_x0y2),
    .MINUS(m2_ch3_aib[75])
   );

  aliasv xaliasv74_ch15 (
    .PLUS(nd_aib74_ch3_x0y2),
    .MINUS(m2_ch3_aib[74])
   );

  aliasv xaliasv73_ch15 (
    .PLUS(nd_aib73_ch3_x0y2),
    .MINUS(m2_ch3_aib[73])
   );

  aliasv xaliasv72_ch15 (
    .PLUS(nd_aib72_ch3_x0y2),
    .MINUS(m2_ch3_aib[72])
   );

  aliasv xaliasv71_ch15 (
    .PLUS(nd_aib71_ch3_x0y2),
    .MINUS(m2_ch3_aib[71])
   );

  aliasv xaliasv70_ch15 (
    .PLUS(nd_aib70_ch3_x0y2),
    .MINUS(m2_ch3_aib[70])
   );

  aliasv xaliasv69_ch15 (
    .PLUS(nd_aib69_ch3_x0y2),
    .MINUS(m2_ch3_aib[69])
   );

  aliasv xaliasv68_ch15 (
    .PLUS(nd_aib68_ch3_x0y2),
    .MINUS(m2_ch3_aib[68])
   );

  aliasv xaliasv67_ch15 (
    .PLUS(nd_aib67_ch3_x0y2),
    .MINUS(m2_ch3_aib[67])
   );

  aliasv xaliasv66_ch15 (
    .PLUS(nd_aib66_ch3_x0y2),
    .MINUS(m2_ch3_aib[66])
   );

  aliasv xaliasv65_ch15 (
    .PLUS(nd_aib65_ch3_x0y2),
    .MINUS(m2_ch3_aib[65])
   );

  aliasv xaliasv64_ch15 (
    .PLUS(nd_aib64_ch3_x0y2),
    .MINUS(m2_ch3_aib[64])
   );

  aliasv xaliasv63_ch15 (
    .PLUS(nd_aib63_ch3_x0y2),
    .MINUS(m2_ch3_aib[63])
   );

  aliasv xaliasv62_ch15 (
    .PLUS(nd_aib62_ch3_x0y2),
    .MINUS(m2_ch3_aib[62])
   );

  aliasv xaliasv61_ch15 (
    .PLUS(nd_aib61_ch3_x0y2),
    .MINUS(m2_ch3_aib[61])
   );

  aliasv xaliasv60_ch15 (
    .PLUS(nd_aib60_ch3_x0y2),
    .MINUS(m2_ch3_aib[60])
   );

  aliasv xaliasv59_ch15 (
    .PLUS(nd_aib59_ch3_x0y2),
    .MINUS(m2_ch3_aib[59])
   );

  aliasv xaliasv58_ch15 (
    .PLUS(nd_aib58_ch3_x0y2),
    .MINUS(m2_ch3_aib[58])
   );

  aliasv xaliasv57_ch15 (
    .PLUS(nd_aib57_ch3_x0y2),
    .MINUS(m2_ch3_aib[57])
   );

  aliasv xaliasv56_ch15 (
    .PLUS(nd_aib56_ch3_x0y2),
    .MINUS(m2_ch3_aib[56])
   );

  aliasv xaliasv55_ch15 (
    .PLUS(nd_aib55_ch3_x0y2),
    .MINUS(m2_ch3_aib[55])
   );

  aliasv xaliasv54_ch15 (
    .PLUS(nd_aib54_ch3_x0y2),
    .MINUS(m2_ch3_aib[54])
   );

  aliasv xaliasv53_ch15 (
    .PLUS(nd_aib53_ch3_x0y2),
    .MINUS(m2_ch3_aib[53])
   );

  aliasv xaliasv52_ch15 (
    .PLUS(nd_aib52_ch3_x0y2),
    .MINUS(m2_ch3_aib[52])
   );

  aliasv xaliasv51_ch15 (
    .PLUS(nd_aib51_ch3_x0y2),
    .MINUS(m2_ch3_aib[51])
   );

  aliasv xaliasv50_ch15 (
    .PLUS(nd_aib50_ch3_x0y2),
    .MINUS(m2_ch3_aib[50])
   );

  aliasv xaliasv49_ch15 (
    .PLUS(nd_aib49_ch3_x0y2),
    .MINUS(m2_ch3_aib[49])
   );

  aliasv xaliasv48_ch15 (
    .PLUS(nd_aib48_ch3_x0y2),
    .MINUS(m2_ch3_aib[48])
   );

  aliasv xaliasv47_ch15 (
    .PLUS(nd_aib47_ch3_x0y2),
    .MINUS(m2_ch3_aib[47])
   );

  aliasv xaliasv46_ch15 (
    .PLUS(nd_aib46_ch3_x0y2),
    .MINUS(m2_ch3_aib[46])
   );

  aliasv xaliasv45_ch15 (
    .PLUS(nd_aib45_ch3_x0y2),
    .MINUS(m2_ch3_aib[45])
   );

  aliasv xaliasv44_ch15 (
    .PLUS(nd_aib44_ch3_x0y2),
    .MINUS(m2_ch3_aib[44])
   );

  aliasv xaliasv43_ch15 (
    .PLUS(nd_aib43_ch3_x0y2),
    .MINUS(m2_ch3_aib[43])
   );

  aliasv xaliasv42_ch15 (
    .PLUS(nd_aib42_ch3_x0y2),
    .MINUS(m2_ch3_aib[42])
   );

  aliasv xaliasv41_ch15 (
    .PLUS(nd_aib41_ch3_x0y2),
    .MINUS(m2_ch3_aib[41])
   );

  aliasv xaliasv40_ch15 (
    .PLUS(nd_aib40_ch3_x0y2),
    .MINUS(m2_ch3_aib[40])
   );

  aliasv xaliasv39_ch15 (
    .PLUS(nd_aib39_ch3_x0y2),
    .MINUS(m2_ch3_aib[39])
   );

  aliasv xaliasv38_ch15 (
    .PLUS(nd_aib38_ch3_x0y2),
    .MINUS(m2_ch3_aib[38])
   );

  aliasv xaliasv37_ch15 (
    .PLUS(nd_aib37_ch3_x0y2),
    .MINUS(m2_ch3_aib[37])
   );

  aliasv xaliasv36_ch15 (
    .PLUS(nd_aib36_ch3_x0y2),
    .MINUS(m2_ch3_aib[36])
   );

  aliasv xaliasv35_ch15 (
    .PLUS(nd_aib35_ch3_x0y2),
    .MINUS(m2_ch3_aib[35])
   );

  aliasv xaliasv34_ch15 (
    .PLUS(nd_aib34_ch3_x0y2),
    .MINUS(m2_ch3_aib[34])
   );

  aliasv xaliasv33_ch15 (
    .PLUS(nd_aib33_ch3_x0y2),
    .MINUS(m2_ch3_aib[33])
   );

  aliasv xaliasv32_ch15 (
    .PLUS(nd_aib32_ch3_x0y2),
    .MINUS(m2_ch3_aib[32])
   );

  aliasv xaliasv31_ch15 (
    .PLUS(nd_aib31_ch3_x0y2),
    .MINUS(m2_ch3_aib[31])
   );

  aliasv xaliasv30_ch15 (
    .PLUS(nd_aib30_ch3_x0y2),
    .MINUS(m2_ch3_aib[30])
   );

  aliasv xaliasv29_ch15 (
    .PLUS(nd_aib29_ch3_x0y2),
    .MINUS(m2_ch3_aib[29])
   );

  aliasv xaliasv28_ch15 (
    .PLUS(nd_aib28_ch3_x0y2),
    .MINUS(m2_ch3_aib[28])
   );

  aliasv xaliasv27_ch15 (
    .PLUS(nd_aib27_ch3_x0y2),
    .MINUS(m2_ch3_aib[27])
   );

  aliasv xaliasv26_ch15 (
    .PLUS(nd_aib26_ch3_x0y2),
    .MINUS(m2_ch3_aib[26])
   );

  aliasv xaliasv25_ch15 (
    .PLUS(nd_aib25_ch3_x0y2),
    .MINUS(m2_ch3_aib[25])
   );

  aliasv xaliasv24_ch15 (
    .PLUS(nd_aib24_ch3_x0y2),
    .MINUS(m2_ch3_aib[24])
   );

  aliasv xaliasv23_ch15 (
    .PLUS(nd_aib23_ch3_x0y2),
    .MINUS(m2_ch3_aib[23])
   );

  aliasv xaliasv22_ch15 (
    .PLUS(nd_aib22_ch3_x0y2),
    .MINUS(m2_ch3_aib[22])
   );

  aliasv xaliasv21_ch15 (
    .PLUS(nd_aib21_ch3_x0y2),
    .MINUS(m2_ch3_aib[21])
   );

  aliasv xaliasv20_ch15 (
    .PLUS(nd_aib20_ch3_x0y2),
    .MINUS(m2_ch3_aib[20])
   );

  aliasv xaliasv19_ch15 (
    .PLUS(nd_aib19_ch3_x0y2),
    .MINUS(m2_ch3_aib[19])
   );

  aliasv xaliasv18_ch15 (
    .PLUS(nd_aib18_ch3_x0y2),
    .MINUS(m2_ch3_aib[18])
   );

  aliasv xaliasv17_ch15 (
    .PLUS(nd_aib17_ch3_x0y2),
    .MINUS(m2_ch3_aib[17])
   );

  aliasv xaliasv16_ch15 (
    .PLUS(nd_aib16_ch3_x0y2),
    .MINUS(m2_ch3_aib[16])
   );

  aliasv xaliasv15_ch15 (
    .PLUS(nd_aib15_ch3_x0y2),
    .MINUS(m2_ch3_aib[15])
   );

  aliasv xaliasv14_ch15 (
    .PLUS(nd_aib14_ch3_x0y2),
    .MINUS(m2_ch3_aib[14])
   );

  aliasv xaliasv13_ch15 (
    .PLUS(nd_aib13_ch3_x0y2),
    .MINUS(m2_ch3_aib[13])
   );

  aliasv xaliasv12_ch15 (
    .PLUS(nd_aib12_ch3_x0y2),
    .MINUS(m2_ch3_aib[12])
   );

  aliasv xaliasv11_ch15 (
    .PLUS(nd_aib11_ch3_x0y2),
    .MINUS(m2_ch3_aib[11])
   );

  aliasv xaliasv10_ch15 (
    .PLUS(nd_aib10_ch3_x0y2),
    .MINUS(m2_ch3_aib[10])
   );

  aliasv xaliasv9_ch15 (
    .PLUS(nd_aib9_ch3_x0y2),
    .MINUS(m2_ch3_aib[9])
   );

  aliasv xaliasv8_ch15 (
    .PLUS(nd_aib8_ch3_x0y2),
    .MINUS(m2_ch3_aib[8])
   );

  aliasv xaliasv7_ch15 (
    .PLUS(nd_aib7_ch3_x0y2),
    .MINUS(m2_ch3_aib[7])
   );

  aliasv xaliasv6_ch15 (
    .PLUS(nd_aib6_ch3_x0y2),
    .MINUS(m2_ch3_aib[6])
   );

  aliasv xaliasv5_ch15 (
    .PLUS(nd_aib5_ch3_x0y2),
    .MINUS(m2_ch3_aib[5])
   );

  aliasv xaliasv4_ch15 (
    .PLUS(nd_aib4_ch3_x0y2),
    .MINUS(m2_ch3_aib[4])
   );

  aliasv xaliasv3_ch15 (
    .PLUS(nd_aib3_ch3_x0y2),
    .MINUS(m2_ch3_aib[3])
   );

  aliasv xaliasv2_ch15 (
    .PLUS(nd_aib2_ch3_x0y2),
    .MINUS(m2_ch3_aib[2])
   );

  aliasv xaliasv1_ch15 (
    .PLUS(nd_aib1_ch3_x0y2),
    .MINUS(m2_ch3_aib[1])
   );

  aliasv xaliasv0_ch15 (
    .PLUS(nd_aib0_ch3_x0y2),
    .MINUS(m2_ch3_aib[0])
   );

endmodule
