// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. 
// Library - aibnd_lib, Cell - aibnd_rxdatapath_rx, View - schematic
// LAST TIME SAVED: Jul  7 14:09:46 2015
// NETLIST TIME: Jul  8 13:09:51 2015
// `timescale 1ns / 1ns 

module aibnd_rxdatapath_rx ( async_dat_outpclk1_1,
     async_dat_outpdir0_1, idat0_in0_dout_clkp, idat1_in0_dout_clkp,
     idataselb_in0_directout2, idataselb_in0_dout_clkp,
     idataselb_outpclk1_1, idataselb_outpdir0_1,
     idirectout_data_outpdir2_1, idlkin_dist_pinp0,
     ilaunch_clk_in0_dout_clkp, irxen_chain1, irxen_inpclk6,
     irxen_inpdir2, irxen_pinp0, istrbclk_pinp0, itxen_in0_directout2,
     itxen_in0_dout_clkp, itxen_outpclk1_1, itxen_outpdir0_1,
     jtag_clkdr_inpclk1n, jtag_clkdr_inpclk6, jtag_clkdr_out_chain1,
     jtag_clkdr_out_diin_clkp, jtag_clkdr_out_directin2,
     jtag_clkdr_out_dirout2, jtag_clkdr_outpclk1_1,
     jtag_clkdr_outpdir0_1, jtag_clkdr_pinp0, jtag_rx_scan_inpclk1n,
     jtag_rx_scan_inpclk6, jtag_rx_scan_out_diin_clkp,
     jtag_rx_scan_out_directin2, jtag_rx_scan_out_dirout2,
     jtag_rx_scan_outpclk1_1, jtag_rx_scan_outpdir0_1,
     jtag_scan_out_chain1, jtag_scan_pinp0, last_bs_out_chain1,
     oclk_inpdir2, oclkb_inpdir2, oclkn_inpdir4, odat0_outpclk1_1,
     odat0_outpdir0_1, odat1_outpclk1_1, odat1_outpdir0_1,
     odat_async_inpclk1, odat_async_inpclk4, odirectin_data,
     odirectin_data_out0_chain1, odll_dll2core_str, odll_lock,
     out_rx_fast_clk, pcs_clk, pcs_data_out0, pcs_data_out1, scan_out,
     shift_en_directout2, shift_en_dout_clkp, shift_en_inpclk1n,
     shift_en_inpclk6, shift_en_inpdir2, shift_en_out_chain1,
     shift_en_outpclk1_1, shift_en_outpdir0_1, shift_en_pinp0,
     iopad_direct_input, iopad_directinclkn, iopad_directinclkp,
     iopad_directout, iopad_directoutclkn, iopad_directoutclkp,
     iopad_inclkn, iopad_inclkp, iopad_indat, avmm_sync_rstb,
     clkdr_xr1l, clkdr_xr1r, clkdr_xr2l, clkdr_xr2r, clkdr_xr3l,
     clkdr_xr3r, clkdr_xr4l, clkdr_xr4r, clkdr_xr5l, clkdr_xr5r,
     clkdr_xr6l, clkdr_xr6r, clkdr_xr7l, clkdr_xr7r, clkdr_xr8l,
     clkdr_xr8r, dft_rx_clk, iasync_dat_outpdir6, iclkin_dist_vinp0,
     iclkin_dist_vinp1, idat0_directoutclkn, idat0_directoutclkp,
     idat0_poutp18, idat1_directoutclkn, idat1_directoutclkp,
     idat1_poutp18, idataselb, idataselb_outpdir6, idataselb_poutp18,
     idatdll_entest_str, idatdll_pipeline_global_en,
     idatdll_rb_clkdiv_str, idatdll_rb_half_code_str,
     idatdll_rb_selflock_str, idatdll_scan_clk_in, idatdll_scan_in,
     idatdll_scan_mode_n, idatdll_scan_rst_n, idatdll_scan_shift_n,
     idatdll_str_align_dyconfig_ctl_static,
     idatdll_str_align_dyconfig_ctlsel,
     idatdll_str_align_stconfig_core_dn_prgmnvrt,
     idatdll_str_align_stconfig_core_up_prgmnvrt,
     idatdll_str_align_stconfig_core_updnen,
     idatdll_str_align_stconfig_dftmuxsel,
     idatdll_str_align_stconfig_dll_en,
     idatdll_str_align_stconfig_dll_rst_en,
     idatdll_str_align_stconfig_hps_ctrl_en,
     idatdll_str_align_stconfig_ndllrst_prgmnvrt,
     idatdll_str_align_stconfig_new_dll,
     idatdll_str_align_stconfig_spare, idatdll_test_clk_pll_en_n,
     iddren_poutp18, idirectout_data, idll_core2dll_str, idll_lock_req,
     ilaunch_clk_poutp18, indrv_r12, indrv_r34, indrv_r56, indrv_r78,
     input_rstb, ipdrv_r12, ipdrv_r34, ipdrv_r56, ipdrv_r78,
     irxen_in_chain1, irxen_inpclk3, irxen_inpdir3, irxen_inpshared0,
     irxen_r0, irxen_r1, irxen_r2, irxen_r3, irxen_vinp0, irxen_vinp1,
     istrbclk_vinp0, istrbclk_vinp1, itxen, itxen_outpdir6,
     itxen_poutp18, jtag_clkdr_in_chain1, jtag_clkdr_inpclk0n,
     jtag_clkdr_inpshared0, jtag_clkdr_out_inpclk3,
     jtag_clkdr_out_inpdir3, jtag_clkdr_out_outpdir6,
     jtag_clkdr_out_poutp18, jtag_clkdr_vinp0, jtag_clkdr_vinp1,
     jtag_clksel, jtag_intest, jtag_mode_in, jtag_rstb, jtag_rstb_en,
     jtag_rx_scan_inpclk0n, jtag_rx_scan_inpshared0,
     jtag_rx_scan_out_inpclk3, jtag_rx_scan_out_inpdir3,
     jtag_rx_scan_out_outpdir6, jtag_rx_scan_out_poutp18,
     jtag_rx_scan_vinp0, jtag_rx_scan_vinp1, jtag_scan_in_chain1,
     jtag_tx_scanen_in, jtag_weakpdn, jtag_weakpu, oclk_inpclk3,
     oclkb_inpclk3, oclkn_inpclk3, oclkn_outpdir4_1, odat0_inpdir0,
     odat1_inpdir0, odat_async_oshared1, odat_async_poutp0,
     odirectin_data_in_chain1, poutp_dig_rstb, rx_shift_en,
     shift_en_in_chain1, shift_en_inpclk0n, shift_en_inpclk3,
     shift_en_inpdir3, shift_en_inpshared0, shift_en_outpdir6,
     shift_en_poutp18, shift_en_vinp0, shift_en_vinp1,
     txdirclk_fast_clkn, txdirclk_fast_clkp, txpma_dig_rstb,
     vccl_aibnd, vssl_aibnd );

output  async_dat_outpclk1_1, async_dat_outpdir0_1,
     idat0_in0_dout_clkp, idat1_in0_dout_clkp,
     idataselb_in0_directout2, idataselb_in0_dout_clkp,
     idataselb_outpclk1_1, idataselb_outpdir0_1,
     idirectout_data_outpdir2_1, idlkin_dist_pinp0,
     ilaunch_clk_in0_dout_clkp, istrbclk_pinp0, itxen_in0_directout2,
     itxen_in0_dout_clkp, itxen_outpclk1_1, itxen_outpdir0_1,
     jtag_clkdr_inpclk1n, jtag_clkdr_inpclk6, jtag_clkdr_out_chain1,
     jtag_clkdr_out_diin_clkp, jtag_clkdr_out_directin2,
     jtag_clkdr_out_dirout2, jtag_clkdr_outpclk1_1,
     jtag_clkdr_outpdir0_1, jtag_clkdr_pinp0, jtag_rx_scan_inpclk1n,
     jtag_rx_scan_inpclk6, jtag_rx_scan_out_diin_clkp,
     jtag_rx_scan_out_directin2, jtag_rx_scan_out_dirout2,
     jtag_rx_scan_outpclk1_1, jtag_rx_scan_outpdir0_1,
     jtag_scan_out_chain1, jtag_scan_pinp0, last_bs_out_chain1,
     oclk_inpdir2, oclkb_inpdir2, oclkn_inpdir4, odat0_outpclk1_1,
     odat0_outpdir0_1, odat1_outpclk1_1, odat1_outpdir0_1,
     odat_async_inpclk1, odat_async_inpclk4,
     odirectin_data_out0_chain1, odll_lock, out_rx_fast_clk, pcs_clk,
     scan_out, shift_en_directout2, shift_en_dout_clkp,
     shift_en_inpclk1n, shift_en_inpclk6, shift_en_inpdir2,
     shift_en_out_chain1, shift_en_outpclk1_1, shift_en_outpdir0_1,
     shift_en_pinp0;

inout  iopad_directinclkn, iopad_directinclkp, iopad_directoutclkn,
     iopad_directoutclkp, iopad_inclkn, iopad_inclkp;

input  avmm_sync_rstb, clkdr_xr1l, clkdr_xr1r, clkdr_xr2l, clkdr_xr2r,
     clkdr_xr3l, clkdr_xr3r, clkdr_xr4l, clkdr_xr4r, clkdr_xr5l,
     clkdr_xr5r, clkdr_xr6l, clkdr_xr6r, clkdr_xr7l, clkdr_xr7r,
     clkdr_xr8l, clkdr_xr8r, dft_rx_clk, iasync_dat_outpdir6,
     iclkin_dist_vinp0, iclkin_dist_vinp1, idat0_directoutclkn,
     idat0_directoutclkp, idat0_poutp18, idat1_directoutclkn,
     idat1_directoutclkp, idat1_poutp18, idataselb_outpdir6,
     idataselb_poutp18, idatdll_entest_str, idatdll_pipeline_global_en,
     idatdll_rb_half_code_str, idatdll_rb_selflock_str,
     idatdll_scan_clk_in, idatdll_scan_in, idatdll_scan_mode_n,
     idatdll_scan_rst_n, idatdll_scan_shift_n,
     idatdll_str_align_dyconfig_ctlsel,
     idatdll_str_align_stconfig_core_dn_prgmnvrt,
     idatdll_str_align_stconfig_core_up_prgmnvrt,
     idatdll_str_align_stconfig_core_updnen,
     idatdll_str_align_stconfig_dll_en,
     idatdll_str_align_stconfig_dll_rst_en,
     idatdll_str_align_stconfig_hps_ctrl_en,
     idatdll_str_align_stconfig_ndllrst_prgmnvrt,
     idatdll_test_clk_pll_en_n, iddren_poutp18, idll_lock_req,
     ilaunch_clk_poutp18, input_rstb, istrbclk_vinp0, istrbclk_vinp1,
     itxen_outpdir6, itxen_poutp18, jtag_clkdr_in_chain1,
     jtag_clkdr_inpclk0n, jtag_clkdr_inpshared0,
     jtag_clkdr_out_inpclk3, jtag_clkdr_out_inpdir3,
     jtag_clkdr_out_outpdir6, jtag_clkdr_out_poutp18, jtag_clkdr_vinp0,
     jtag_clkdr_vinp1, jtag_clksel, jtag_intest, jtag_mode_in,
     jtag_rstb, jtag_rstb_en, jtag_rx_scan_inpclk0n,
     jtag_rx_scan_inpshared0, jtag_rx_scan_out_inpclk3,
     jtag_rx_scan_out_inpdir3, jtag_rx_scan_out_outpdir6,
     jtag_rx_scan_out_poutp18, jtag_rx_scan_vinp0, jtag_rx_scan_vinp1,
     jtag_scan_in_chain1, jtag_tx_scanen_in, jtag_weakpdn, jtag_weakpu,
     oclk_inpclk3, oclkb_inpclk3, oclkn_inpclk3, oclkn_outpdir4_1,
     odat0_inpdir0, odat1_inpdir0, odat_async_oshared1,
     odat_async_poutp0, odirectin_data_in_chain1, poutp_dig_rstb,
     shift_en_in_chain1, shift_en_inpclk0n, shift_en_inpclk3,
     shift_en_inpdir3, shift_en_inpshared0, shift_en_outpdir6,
     shift_en_poutp18, shift_en_vinp0, shift_en_vinp1,
     txdirclk_fast_clkn, txdirclk_fast_clkp, txpma_dig_rstb,
     vccl_aibnd, vssl_aibnd;

output [2:0]  irxen_pinp0;
output [2:0]  irxen_inpclk6;
output [2:0]  irxen_inpdir2;
output [2:0]  irxen_chain1;
output [12:0]  odll_dll2core_str;
output [6:0]  odirectin_data;
output [19:0]  pcs_data_out1;
output [19:0]  pcs_data_out0;

inout [19:0]  iopad_indat;
inout [3:0]  iopad_directout;
inout [6:0]  iopad_direct_input;

input [2:0]  idll_core2dll_str;
input [2:0]  irxen_inpshared0;
input [1:0]  indrv_r34;
input [9:0]  idatdll_str_align_dyconfig_ctl_static;
input [2:0]  idatdll_rb_clkdiv_str;
input [2:0]  irxen_inpclk3;
input [2:0]  irxen_vinp0;
input [1:0]  indrv_r56;
input [1:0]  ipdrv_r56;
input [2:0]  irxen_inpdir3;
input [1:0]  ipdrv_r34;
input [1:0]  ipdrv_r12;
input [2:0]  irxen_r2;
input [2:0]  itxen;
input [3:0]  idirectout_data;
input [1:0]  indrv_r12;
input [2:0]  irxen_r1;
input [10:0]  idatdll_str_align_stconfig_spare;
input [2:0]  irxen_r0;
input [19:0]  idatdll_str_align_stconfig_dftmuxsel;
input [1:0]  ipdrv_r78;
input [1:0]  indrv_r78;
input [2:0]  idataselb;
input [2:0]  irxen_vinp1;
input [2:0]  irxen_in_chain1;
input [2:0]  irxen_r3;
input [2:0]  idatdll_str_align_stconfig_new_dll;
input [36:0]  rx_shift_en;

wire dll_scan_out, scan_out, pcs_clk_inv, lstrbclk_rep ; // Conversion Sript Generated

// Buses in the design

wire  [1:2]  nc_odat0_out0_directout;

wire  [1:1]  nc_oclkn_out0_directin;

wire  [0:1]  nc_oclk_out0_directin;

wire  [0:3]  nc_pd_data_directout;

wire  [1:6]  nc_odata0_out0_directin;

wire  [51:0]  csr_reg_str;

wire  [0:19]  pcs_data_out0_io;

wire  [0:6]  nc_oclk_directin;

wire  [1:2]  nc_odat1_out0_directout;

wire  [12:12]  ncdrx_oclkb;

wire  [12:12]  ncdrx_oclkn;

wire  [12:12]  ncdrx_oclk;

wire  [0:11]  rx_strbclk_l;

wire  [0:1]  odirectin_data_out0;

wire  [0:1]  nc_oclkb_out0_directin;

wire  [0:11]  rx_distclk_l;

wire  [0:6]  nc_pd_data_out0_directin;

wire  [0:6]  nc_odata0_directin;

wire  [0:6]  nc_oclkb_directin;

wire  [0:19]  pcs_data_out1_io;

wire  [0:3]  nc_odat1_directout;

wire  [0:3]  nc_odat_async_directout;

wire  [0:3]  nc_oclk_directout;

wire  [0:3]  nc_oclkb_directout;

wire  [0:3]  nc_pd_data_out0_directout;

wire  [0:11]  rx_strbclk_r;

wire  [1:6]  nc_odata1_out0_directin;

wire  [0:11]  rx_distclk_r;

wire  [0:6]  nc_odata1_directin;

wire  [0:3]  nc_oclkb_out0_directout;

wire  [0:3]  nc_oclk_out0_directout;

wire  [0:3]  nc_odat_async_out0_directout;

wire  [0:6]  nc_pd_data_directin;

wire  [0:3]  nc_odat0_directout;

wire  [0:3]  nc_oclkn_out0_directout;


// specify 
//     specparam CDS_LIBNAME  = "aibnd_lib";
//     specparam CDS_CELLNAME = "aibnd_rxdatapath_rx";
//     specparam CDS_VIEWNAME = "schematic";
// endspecify
wire oclk_clkp_buf;
wire oclk_clkpb_buf;
wire oclk_clkp_io;
wire oclk_clkpb_io;

aibnd_clktree_pcs  clktree_pcs ( /*.vcc_aibnd(vccl_aibnd),
     .vss_aibnd(vssl_aibnd),*/ .lstrbclk_mimic2(clk_distclk),
     .lstrbclk_r_11(rx_distclk_r[11]),
     .lstrbclk_r_10(rx_distclk_r[10]), .lstrbclk_r_9(rx_distclk_r[9]),
     .lstrbclk_r_8(rx_distclk_r[8]), .lstrbclk_r_7(rx_distclk_r[7]),
     .lstrbclk_r_6(rx_distclk_r[6]), .lstrbclk_r_5(rx_distclk_r[5]),
     .lstrbclk_r_4(rx_distclk_r[4]), .lstrbclk_r_3(rx_distclk_r[3]),
     .lstrbclk_r_2(rx_distclk_r[2]), .lstrbclk_r_1(rx_distclk_r[1]),
     .lstrbclk_r_0(rx_distclk_r[0]), .lstrbclk_mimic1(nc_clk_mimic1),
     .lstrbclk_mimic0(nc_clk_mimic0), .lstrbclk_l_0(rx_distclk_l[0]),
     .lstrbclk_l_1(rx_distclk_l[1]), .lstrbclk_l_2(rx_distclk_l[2]),
     .lstrbclk_l_3(rx_distclk_l[3]), .lstrbclk_l_4(rx_distclk_l[4]),
     .lstrbclk_l_5(rx_distclk_l[5]), .lstrbclk_l_6(rx_distclk_l[6]),
     .lstrbclk_l_7(rx_distclk_l[7]), .lstrbclk_l_8(rx_distclk_l[8]),
     .lstrbclk_l_9(rx_distclk_l[9]), .lstrbclk_l_10(rx_distclk_l[10]),
     .lstrbclk_l_11(rx_distclk_l[11]), .lstrbclk_rep(lstrbclk_rep),
     .clkin(oclk_clkp_buf));
aibnd_aliasd  aliasd11 ( .MINUS(shift_en_inpclk6), .PLUS(rx_shift_en[3]));
aibnd_aliasd  aliasv99[2:0] ( .MINUS(irxen_chain1[2:0]),      .PLUS(irxen_r2[2:0]));
aibnd_aliasd  aliasd4 ( .MINUS(shift_en_pinp0), .PLUS(rx_shift_en[33]));
aibnd_aliasd  aliasd10 ( .MINUS(shift_en_inpclk1n), .PLUS(rx_shift_en[8]));
aibnd_aliasd  aliasv55 ( .MINUS(idataselb_in0_directout2),      .PLUS(idataselb[1]));
aibnd_aliasd  aliasd3[2:0] ( .MINUS(irxen_inpclk6[2:0]),      .PLUS(irxen_r2[2:0]));
aibnd_aliasd  aliasd1[2:0] ( .MINUS(irxen_pinp0[2:0]), .PLUS(irxen_r0[2:0]));
aibnd_aliasd  aliasd2 ( .MINUS(istrbclk_pinp0),      .PLUS(rx_strbclk_r[11]));
aibnd_aliasd  aliasv41 ( .MINUS(itxen_in0_dout_clkp), .PLUS(itxen[0]));
aibnd_aliasd  aliasd0 ( .MINUS(idlkin_dist_pinp0),      .PLUS(rx_distclk_r[11]));
aibnd_aliasd  aliasv88 ( .MINUS(csr_reg_str[51]),      .PLUS(idatdll_str_align_stconfig_hps_ctrl_en));
aibnd_aliasd  aliasv86 ( .MINUS(csr_reg_str[1]),      .PLUS(idatdll_str_align_stconfig_dll_en));
aibnd_aliasd  aliasv85[2:0] ( .MINUS(csr_reg_str[50:48]),      .PLUS(idatdll_str_align_stconfig_new_dll[2:0]));
aibnd_aliasd  aliasv87 ( .MINUS(csr_reg_str[0]),      .PLUS(idatdll_str_align_stconfig_dll_rst_en));
aibnd_aliasd  aliasv53 ( .MINUS(itxen_in0_directout2), .PLUS(itxen[1]));
aibnd_aliasd  aliasv37 ( .MINUS(ilaunch_clk_in0_dout_clkp),      .PLUS(txdirclk_fast_clkp));
aibnd_aliasd  aliasd5 ( .MINUS(shift_en_out_chain1), .PLUS(rx_shift_en[36]));
aibnd_aliasd  aliasv28[2:0] ( .MINUS(irxen_inpdir2[2:0]),      .PLUS(irxen_r2[2:0]));
aibnd_aliasd  aliasd6 ( .MINUS(shift_en_directout2), .PLUS(rx_shift_en[9]));
aibnd_aliasd  aliasv30 ( .MINUS(idataselb_outpclk1_1), .PLUS(idataselb[1]));
aibnd_aliasd  aliasd7 ( .MINUS(shift_en_dout_clkp), .PLUS(rx_shift_en[4]));
aibnd_aliasd  aliasd8 ( .MINUS(shift_en_outpdir0_1), .PLUS(rx_shift_en[11]));
aibnd_aliasd  aliasv96[9:0] ( .MINUS(csr_reg_str[27:18]),      .PLUS(idatdll_str_align_dyconfig_ctl_static[9:0]));
aibnd_aliasd  aliasv95 ( .MINUS(csr_reg_str[17]),      .PLUS(idatdll_str_align_dyconfig_ctlsel));
aibnd_aliasd  aliasv94[10:0] ( .MINUS(csr_reg_str[16:6]),      .PLUS(idatdll_str_align_stconfig_spare[10:0]));
aibnd_aliasd  aliasv93 ( .MINUS(csr_reg_str[5]),      .PLUS(idatdll_str_align_stconfig_core_updnen));
aibnd_aliasd  aliasv92 ( .MINUS(csr_reg_str[4]),      .PLUS(idatdll_str_align_stconfig_core_dn_prgmnvrt));
aibnd_aliasd  aliasv91 ( .MINUS(csr_reg_str[3]),      .PLUS(idatdll_str_align_stconfig_core_up_prgmnvrt));
aibnd_aliasd  aliasd12 ( .MINUS(shift_en_inpdir2), .PLUS(rx_shift_en[0]));
aibnd_aliasd  aliasv71 ( .MINUS(idataselb_outpdir0_1), .PLUS(idataselb[1]));
aibnd_aliasd  aliasv66 ( .MINUS(itxen_outpdir0_1), .PLUS(itxen[1]));
aibnd_aliasd  aliasv36 ( .MINUS(idataselb_in0_dout_clkp),      .PLUS(idataselb[0]));
aibnd_aliasd  aliasv89[19:0] ( .MINUS(csr_reg_str[47:28]),      .PLUS(idatdll_str_align_stconfig_dftmuxsel[19:0]));
aibnd_aliasd  aliasv90 ( .MINUS(csr_reg_str[2]),      .PLUS(idatdll_str_align_stconfig_ndllrst_prgmnvrt));
aibnd_aliasd  aliasv35 ( .MINUS(itxen_outpclk1_1), .PLUS(itxen[1]));
aibnd_aliasd  aliasd9 ( .MINUS(shift_en_outpclk1_1), .PLUS(rx_shift_en[10]));
aibnd_buffx1_top xdirect_in6 ( .idata1_in1_jtag_out(nc_idat1_inpclk2),
     .async_dat_in1_jtag_out(nc_async_dat_inpclk2),
     .idata0_in1_jtag_out(nc_idat0_inpclk2),
     .jtag_clkdr_outn(jtag_clkdr_outn_inpclk2),
     .prev_io_shift_en(rx_shift_en[7]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_directin[6]),
     .oclk_out(nc_oclk_directin[6]), .oclkb_out(nc_oclkb_directin[6]),
     .odat0_out(nc_odata0_directin[6]),
     .odat1_out(nc_odata1_directin[6]),
     .odat_async_out(odirectin_data[6]),
     .pd_data_out(nc_pd_data_directin[6]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(vssl_aibnd),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vssl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r2[2:0]), .irxen_in1(irxen_r3[2:0]),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odata_async_out0_directin6),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(odat_async_inpclk5),
     .shift_en(rx_shift_en[1]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(input_rstb), .jtag_clkdr_out(jtag_clkdr_out_inpclk2),
     .odat1_aib(nc_odata1_out0_directin[6]),
     .jtag_rx_scan_out(jtag_rx_scan_out_inpclk2),
     .odat0_aib(nc_odata0_out0_directin[6]),
     .oclk_aib(oclk_out0_directin6),
     .last_bs_out(nc_last_bs_out_inpclk2),
     .oclkb_aib(oclkb_out0_directin6), .jtag_clkdr_in(clkdr_xr1l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_inpclk1),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_direct_input[6]), .oclkn(nc_oclkn_out0_directin6),
     .iclkn(oclkn_inpclk3), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdirect_out3 (
     .idata1_in1_jtag_out(nc_idat1_outpdir0_1),
     .async_dat_in1_jtag_out(async_dat_outpdir0_1),
     .idata0_in1_jtag_out(nc_idat0_outpdir0_1),
     .jtag_clkdr_outn(jtag_clkdr_outn_outpdir0_1),
     .prev_io_shift_en(shift_en_vinp1), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb),
     .pd_data_aib(nc_pd_data_out0_directout[3]),
     .oclk_out(nc_oclk_directout[3]),
     .oclkb_out(nc_oclkb_directout[3]),
     .odat0_out(nc_odat0_directout[3]),
     .odat1_out(nc_odat1_directout[3]),
     .odat_async_out(nc_odat_async_directout[3]),
     .pd_data_out(nc_pd_data_directout[3]),
     .async_dat_in0(idirectout_data[3]), .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(iclkin_dist_vinp1),
     .iclkin_dist_in1(iclkin_dist_vinp1), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(idataselb[1]),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r12[1:0]),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0(ipdrv_r12[1:0]),
     .ipdrv_in1({vssl_aibnd, vssl_aibnd}), .irxen_in0({vssl_aibnd,
     vccl_aibnd, vssl_aibnd}), .irxen_in1(irxen_vinp1[2:0]),
     .istrbclk_in0(istrbclk_vinp1), .istrbclk_in1(istrbclk_vinp1),
     .itxen_in0(itxen[1]), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_out0_directout[3]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[11]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(avmm_sync_rstb), .jtag_clkdr_out(jtag_clkdr_outpdir0_1),
     .odat1_aib(odat1_outpdir0_1),
     .jtag_rx_scan_out(jtag_rx_scan_outpdir0_1),
     .odat0_aib(odat0_outpdir0_1),
     .oclk_aib(nc_oclk_out0_directout[3]),
     .last_bs_out(nc_last_bs_out_directout3),
     .oclkb_aib(nc_oclkb_out0_directout[3]),
     .jtag_clkdr_in(clkdr_xr2l), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_vinp1),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_directout[3]), .oclkn(nc_oclkn_out0_directout[3]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdirect_out1 (
     .idata1_in1_jtag_out(nc_idat1_directout1),
     .async_dat_in1_jtag_out(async_dat_directout1),
     .idata0_in1_jtag_out(nc_idat0_directout1),
     .jtag_clkdr_outn(jtag_clkdr_outn_directout1),
     .prev_io_shift_en(shift_en_poutp18), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb),
     .pd_data_aib(nc_pd_data_out0_directout[1]),
     .oclk_out(nc_oclk_directout[1]),
     .oclkb_out(nc_oclkb_directout[1]),
     .odat0_out(nc_odat0_directout[1]),
     .odat1_out(nc_odat1_directout[1]),
     .odat_async_out(nc_odat_async_directout[1]),
     .pd_data_out(nc_pd_data_directout[1]),
     .async_dat_in0(idirectout_data[1]), .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(vssl_aibnd), .iclkin_dist_in1(vssl_aibnd),
     .idata0_in0(vssl_aibnd), .idata0_in1(idat0_poutp18),
     .idata1_in0(vssl_aibnd), .idata1_in1(idat1_poutp18),
     .idataselb_in0(idataselb[1]), .idataselb_in1(idataselb_poutp18),
     .iddren_in0(vssl_aibnd), .iddren_in1(iddren_poutp18),
     .ilaunch_clk_in0(ilaunch_clk_poutp18),
     .ilaunch_clk_in1(ilaunch_clk_poutp18), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r56[1:0]),
     .indrv_in1(indrv_r56[1:0]), .ipdrv_in0(ipdrv_r56[1:0]),
     .ipdrv_in1(ipdrv_r56[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[1]), .itxen_in1(itxen_poutp18),
     .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_out0_directout[1]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[12]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(txpma_dig_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_directout1),
     .odat1_aib(nc_odat1_out0_directout[1]),
     .jtag_rx_scan_out(jtag_rx_scan_out_directout1),
     .odat0_aib(nc_odat0_out0_directout[1]),
     .oclk_aib(nc_oclk_out0_directout[1]),
     .last_bs_out(nc_last_bs_out_directout1),
     .oclkb_aib(nc_oclkb_out0_directout[1]),
     .jtag_clkdr_in(clkdr_xr5l), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_poutp18),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_directout[1]), .oclkn(nc_oclkn_out0_directout[1]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp0 ( .idata1_in1_jtag_out(nc_idat1_pinp0),
     .async_dat_in1_jtag_out(nc_async_dat_pinp0),
     .idata0_in1_jtag_out(nc_idat0_pinp0),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp0),
     .prev_io_shift_en(rx_shift_en[31]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(pd_data__out0_pinp0),
     .oclk_out(nc_oclk_pinp0), .oclkb_out(nc_oclkb_pinp0),
     .odat0_out(pcs_data_out0_io[0]), .odat1_out(pcs_data_out1_io[0]),
     .odat_async_out(nc_odat_async_pinp0),
     .pd_data_out(nc_pd_data_pinp0), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_r[7]),
     .iclkin_dist_in1(rx_distclk_r[7]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(rx_strbclk_r[7]), .istrbclk_in1(rx_strbclk_r[7]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(odirectin_data_out0_pinp0),
     .oclkb_in1(vssl_aibnd), .odat0_in1(odat0_inpdir0),
     .odat1_in1(odat1_inpdir0), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[33]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_pinp0),
     .odat1_aib(ncdrx_odat1_out0_pinp0),
     .jtag_rx_scan_out(jtag_scan_pinp0),
     .odat0_aib(ncdrx_odat0_out0_pinp0),
     .oclk_aib(ncdrx_oclk_out0_pinp0), .last_bs_out(last_bs_out_pinp0),
     .oclkb_aib(ncdrx_oclkb_out0_pinp0), .jtag_clkdr_in(clkdr_xr7r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_pinp2),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp2), .iopad(iopad_indat[0]),
     .oclkn(ncdrx_oclkn_out0_pinp0), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp2 ( .idata1_in1_jtag_out(nc_idat1_pinp2),
     .async_dat_in1_jtag_out(nc_async_dat_pinp2),
     .idata0_in1_jtag_out(nc_idat0_pinp2),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp2),
     .prev_io_shift_en(rx_shift_en[29]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(pd_data__out0_pinp2),
     .oclk_out(nc_oclk_pinp2), .oclkb_out(nc_oclkb_pinp2),
     .odat0_out(pcs_data_out0_io[2]), .odat1_out(pcs_data_out1_io[2]),
     .odat_async_out(nc_odat_async_pinp2),
     .pd_data_out(nc_pd_data_pinp2), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_r[3]),
     .iclkin_dist_in1(rx_distclk_r[3]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(rx_strbclk_r[3]), .istrbclk_in1(rx_strbclk_r[3]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(odirectin_data_out0_pinp2),
     .oclkb_in1(vssl_aibnd), .odat0_in1(ncdrx_odat0_out0_pinp0),
     .odat1_in1(ncdrx_odat1_out0_pinp0), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[31]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_pinp2),
     .odat1_aib(ncdrx_odat1_out0_pinp2),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp2),
     .odat0_aib(ncdrx_odat0_out0_pinp2),
     .oclk_aib(ncdrx_oclk_out0_pinp2), .last_bs_out(last_bs_out_pinp2),
     .oclkb_aib(ncdrx_oclkb_out0_pinp2), .jtag_clkdr_in(clkdr_xr7r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_pinp4),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp4), .iopad(iopad_indat[2]),
     .oclkn(ncdrx_oclkn_out0_pinp2), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp4 ( .idata1_in1_jtag_out(nc_idat1_pinp4),
     .async_dat_in1_jtag_out(nc_async_dat_pinp4),
     .idata0_in1_jtag_out(nc_idat0_pinp4),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp4),
     .prev_io_shift_en(rx_shift_en[27]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_pinp4),
     .oclk_out(nc_oclk_pinp4), .oclkb_out(nc_oclkb_pinp4),
     .odat0_out(pcs_data_out0_io[4]), .odat1_out(pcs_data_out1_io[4]),
     .odat_async_out(nc_odat_async_pinp4),
     .pd_data_out(nc_pd_data_pinp4), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_r[1]),
     .iclkin_dist_in1(rx_distclk_r[1]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(rx_strbclk_r[1]), .istrbclk_in1(rx_strbclk_r[1]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(nc_odat_async_out0_pinp4),
     .oclkb_in1(vssl_aibnd), .odat0_in1(ncdrx_odat0_out0_pinp2),
     .odat1_in1(ncdrx_odat1_out0_pinp2), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[29]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_pinp4),
     .odat1_aib(ncdrx_odat1_pinp4),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp4),
     .odat0_aib(ncdrx_odat0_pinp4), .oclk_aib(ncdrx_oclk_pinp4),
     .last_bs_out(last_bs_out_pinp4), .oclkb_aib(ncdrx_oclkb_pinp4),
     .jtag_clkdr_in(clkdr_xr7r), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_pinp6),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp6), .iopad(iopad_indat[4]),
     .oclkn(ncdrx_oclkn_pinp4), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp6 ( .idata1_in1_jtag_out(nc_idat1_pinp6),
     .async_dat_in1_jtag_out(nc_async_dat_pinp6),
     .idata0_in1_jtag_out(nc_idat0_pinp6),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp6),
     .prev_io_shift_en(rx_shift_en[25]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_pinp6),
     .oclk_out(nc_oclk_pinp6), .oclkb_out(nc_oclkb_pinp6),
     .odat0_out(pcs_data_out0_io[6]), .odat1_out(pcs_data_out1_io[6]),
     .odat_async_out(nc_odat_async_pinp6),
     .pd_data_out(nc_pd_data_pinp6), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_r[5]),
     .iclkin_dist_in1(rx_distclk_r[5]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(rx_strbclk_r[5]), .istrbclk_in1(rx_strbclk_r[5]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(nc_odat_async_out0_pinp6),
     .oclkb_in1(vssl_aibnd), .odat0_in1(ncdrx_odat0_pinp4),
     .odat1_in1(ncdrx_odat1_pinp4), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[27]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_pinp6),
     .odat1_aib(pcs_data_out1_pinp6),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp6),
     .odat0_aib(pcs_data_out0_pinp6), .oclk_aib(nc_oclk_out0_pinp6),
     .last_bs_out(last_bs_out_pinp6), .oclkb_aib(nc_oclkb_out0_pinp6),
     .jtag_clkdr_in(clkdr_xr7r), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_pinp8),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp8), .iopad(iopad_indat[6]),
     .oclkn(nc_oclkn_out0_pinp6), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp8 ( .idata1_in1_jtag_out(nc_idat1_pinp8),
     .async_dat_in1_jtag_out(nc_async_dat_pinp8),
     .idata0_in1_jtag_out(nc_idat0_pinp8),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp8),
     .prev_io_shift_en(rx_shift_en[23]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_pinp8),
     .oclk_out(nc_oclk_pinp8), .oclkb_out(nc_oclkb_pinp8),
     .odat0_out(pcs_data_out0_io[8]), .odat1_out(pcs_data_out1_io[8]),
     .odat_async_out(nc_odat_async_pinp8),
     .pd_data_out(nc_pd_data_pinp8), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_r[9]),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(idat0_rx_clkp), .idata1_in0(vssl_aibnd),
     .idata1_in1(idat1_rx_clkp), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vccl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vccl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(dft_rx_clk), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1(irxen_r1[2:0]),
     .istrbclk_in0(rx_strbclk_r[9]), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(nc_odat_async_out0_pinp8),
     .oclkb_in1(vssl_aibnd), .odat0_in1(pcs_data_out0_pinp6),
     .odat1_in1(pcs_data_out1_pinp6), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[25]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_pinp8),
     .odat1_aib(ncdrx_odat1_pinp8),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp8),
     .odat0_aib(ncdrx_odat0_pinp8), .oclk_aib(oclk_pinp8),
     .last_bs_out(last_bs_out_pinp8), .oclkb_aib(oclkb_pinp8),
     .jtag_clkdr_in(clkdr_xr7r), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(nc_jtag_rx_scan_out_rx_clkp),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(nc_last_bs_out_rx_clkp), .iopad(iopad_indat[8]),
     .oclkn(ncdrx_oclkn_pinp8), .iclkn(oclkn_pinp9),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xrx_clkp ( .idata1_in1_jtag_out(idat1_rx_clkp),
     .async_dat_in1_jtag_out(nc_async_dat_rx_clkp),
     .idata0_in1_jtag_out(idat0_rx_clkp),
     .jtag_clkdr_outn(jtag_clkdr_outn_rx_clkp),
     .prev_io_shift_en(rx_shift_en[21]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(pd_data_out0_rx_clkp),
     .oclk_out(oclk_clkp_io), .oclkb_out(oclk_clkpb_io),
     .odat0_out(nc_odat0_rx_clkp), .odat1_out(nc_odat1__rx_clkp),
     .odat_async_out(nc_odat_async_rx_clkp),
     .pd_data_out(nc_pd_data_rx_clkp), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_l[11]),
     .iclkin_dist_in1(rx_distclk_l[11]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vccl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(dft_rx_clk),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r1[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(rx_strbclk_l[11]), .istrbclk_in1(rx_strbclk_l[11]),
     .itxen_in0(idatdll_str_align_stconfig_spare[0]),
     .itxen_in1(vssl_aibnd), .oclk_in1(oclk_clkp_buf),
     .odat_async_aib(ncdrx_odat_async_out0_rx_clkp),
     .oclkb_in1(oclk_clkpb_buf), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[23]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb),
     .jtag_clkdr_out(nc_jtag_clkdr_out_rx_clkp),
     .odat1_aib(drx_odat1_out0_rx_clkp),
     .jtag_rx_scan_out(nc_jtag_rx_scan_out_rx_clkp),
     .odat0_aib(drx_odat0_out0_rx_clkp),
     .oclk_aib(drx_oclk_out0_rx_clkp),
     .last_bs_out(nc_last_bs_out_rx_clkp),
     .oclkb_aib(drx_oclkb_out0_rx_clkp), .jtag_clkdr_in(clkdr_xr7l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_pinp10),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp10), .iopad(iopad_inclkp),
     .oclkn(ncdrx_oclkn_rx_clkp), .iclkn(oclkn_clkn),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp10 ( .idata1_in1_jtag_out(nc_idat1_pinp10),
     .async_dat_in1_jtag_out(nc_async_dat_pinp10),
     .idata0_in1_jtag_out(nc_idat0_pinp10),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp10),
     .prev_io_shift_en(rx_shift_en[19]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(pd_data__out0_pinp10),
     .oclk_out(nc_oclk_pinp10), .oclkb_out(nc_oclkb_pinp10),
     .odat0_out(pcs_data_out0_io[10]),
     .odat1_out(pcs_data_out1_io[10]),
     .odat_async_out(nc_odat_async_pinp10),
     .pd_data_out(nc_pd_data_pinp10), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_l[7]),
     .iclkin_dist_in1(rx_distclk_l[7]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(rx_strbclk_l[7]), .istrbclk_in1(rx_strbclk_l[7]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd),
     .odat_async_aib(odirectin_data_out0_pinp10),
     .oclkb_in1(vssl_aibnd), .odat0_in1(drx_odat0_out0_rx_clkp),
     .odat1_in1(drx_odat1_out0_rx_clkp), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[21]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_pinp10),
     .odat1_aib(odat1_pinp10),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp10),
     .odat0_aib(odat0_pinp10), .oclk_aib(ncdrx_oclk_out0_pinp10),
     .last_bs_out(last_bs_out_pinp10),
     .oclkb_aib(ncdrx_oclkb_out0_pinp10), .jtag_clkdr_in(clkdr_xr7l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_pinp12),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp12), .iopad(iopad_indat[10]),
     .oclkn(ncdrx_oclkn_out0_pinp10), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp12 ( .idata1_in1_jtag_out(nc_idat1_pinp12),
     .async_dat_in1_jtag_out(nc_async_dat_pinp12),
     .idata0_in1_jtag_out(nc_idat0_pinp12),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp12),
     .prev_io_shift_en(rx_shift_en[17]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(pd_data__out0_pinp12),
     .oclk_out(nc_oclk_pinp12), .oclkb_out(nc_oclkb_pinp12),
     .odat0_out(pcs_data_out0_io[12]),
     .odat1_out(pcs_data_out1_io[12]),
     .odat_async_out(nc_odat_async_pinp12),
     .pd_data_out(nc_pd_data_pinp12), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_l[3]),
     .iclkin_dist_in1(rx_distclk_l[3]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(rx_strbclk_l[3]), .istrbclk_in1(rx_strbclk_l[3]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd),
     .odat_async_aib(odirectin_data_out0_pinp12),
     .oclkb_in1(vssl_aibnd), .odat0_in1(odat0_pinp10),
     .odat1_in1(odat1_pinp10), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[19]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_pinp12),
     .odat1_aib(odat1_pinp12),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp12),
     .odat0_aib(odat0_pinp12), .oclk_aib(ncdrx_oclk[12]),
     .last_bs_out(last_bs_out_pinp12), .oclkb_aib(ncdrx_oclkb[12]),
     .jtag_clkdr_in(clkdr_xr7l), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_pinp14),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp14), .iopad(iopad_indat[12]),
     .oclkn(ncdrx_oclkn[12]), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp14 ( .idata1_in1_jtag_out(nc_idat1_pinp14),
     .async_dat_in1_jtag_out(nc_async_dat_pinp14),
     .idata0_in1_jtag_out(nc_idat0_pinp14),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp14),
     .prev_io_shift_en(rx_shift_en[15]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(pd_data__out0_pinp14),
     .oclk_out(nc_oclk_pinp14), .oclkb_out(nc_oclkb_pinp14),
     .odat0_out(pcs_data_out0_io[14]),
     .odat1_out(pcs_data_out1_io[14]),
     .odat_async_out(nc_odat_async_pinp14),
     .pd_data_out(nc_pd_data_pinp14), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_l[1]),
     .iclkin_dist_in1(rx_distclk_l[1]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(rx_strbclk_l[1]), .istrbclk_in1(rx_strbclk_l[1]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd),
     .odat_async_aib(odirectin_data_out0_pinp14),
     .oclkb_in1(vssl_aibnd), .odat0_in1(odat0_pinp12),
     .odat1_in1(odat1_pinp12), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[17]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_pinp14),
     .odat1_aib(odat1_pinp14),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp14),
     .odat0_aib(odat0_pinp14), .oclk_aib(ncdrx_oclk_pinp14),
     .last_bs_out(last_bs_out_pinp14), .oclkb_aib(ncdrx_oclkb_pinp14),
     .jtag_clkdr_in(clkdr_xr7l), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_pinp16),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp16), .iopad(iopad_indat[14]),
     .oclkn(ncdrx_oclkn_pinp14), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp16 ( .idata1_in1_jtag_out(nc_idat1_pinp16),
     .async_dat_in1_jtag_out(nc_async_dat_pinp16),
     .idata0_in1_jtag_out(nc_idat0_pinp16),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp16),
     .prev_io_shift_en(rx_shift_en[13]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_pinp16),
     .oclk_out(nc_oclk_pinp16), .oclkb_out(nc_oclkb_pinp16),
     .odat0_out(pcs_data_out0_io[16]),
     .odat1_out(pcs_data_out1_io[16]),
     .odat_async_out(nc_odat_async_pinp16),
     .pd_data_out(nc_pd_data_pinp16), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_l[5]),
     .iclkin_dist_in1(rx_distclk_l[5]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(rx_strbclk_l[5]), .istrbclk_in1(rx_strbclk_l[5]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(nc_odat_async_out0_pinp16),
     .oclkb_in1(vssl_aibnd), .odat0_in1(odat0_pinp14),
     .odat1_in1(odat1_pinp14), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[15]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_pinp16),
     .odat1_aib(pcs_data_out1_pinp16),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp16),
     .odat0_aib(pcs_data_out0_pinp16), .oclk_aib(nc_oclk_out0_pinp16),
     .last_bs_out(last_bs_out_pinp16),
     .oclkb_aib(nc_oclkb_out0_pinp16), .jtag_clkdr_in(clkdr_xr7l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_pinp18),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp18), .iopad(iopad_indat[16]),
     .oclkn(nc_oclkn_out0_pinp16), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp18 ( .idata1_in1_jtag_out(nc_idat1_pinp18),
     .async_dat_in1_jtag_out(nc_async_dat_pinp18),
     .idata0_in1_jtag_out(nc_idat0_pinp18),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp18),
     .prev_io_shift_en(rx_shift_en[12]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(pd_data_pinp18),
     .oclk_out(nc_oclk_pinp18), .oclkb_out(nc_oclkb_pinp18),
     .odat0_out(pcs_data_out0_io[18]),
     .odat1_out(pcs_data_out1_io[18]),
     .odat_async_out(nc_odat_async_pinp18),
     .pd_data_out(nc_pd_data_pinp18), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(async_dat_directout1),
     .iclkin_dist_in0(rx_distclk_l[9]), .iclkin_dist_in1(vssl_aibnd),
     .idata0_in0(vssl_aibnd), .idata0_in1(vssl_aibnd),
     .idata1_in0(vssl_aibnd), .idata1_in1(vssl_aibnd),
     .idataselb_in0(vccl_aibnd), .idataselb_in1(idataselb[1]),
     .iddren_in0(vccl_aibnd), .iddren_in1(vssl_aibnd),
     .ilaunch_clk_in0(vssl_aibnd), .ilaunch_clk_in1(vssl_aibnd),
     .ilpbk_dat_in0(vssl_aibnd), .ilpbk_dat_in1(vssl_aibnd),
     .ilpbk_en_in0(vssl_aibnd), .ilpbk_en_in1(vssl_aibnd),
     .indrv_in0({vssl_aibnd, vssl_aibnd}), .indrv_in1(indrv_r78[1:0]),
     .ipdrv_in0({vssl_aibnd, vssl_aibnd}), .ipdrv_in1(ipdrv_r78[1:0]),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .istrbclk_in0(rx_strbclk_l[9]),
     .istrbclk_in1(vssl_aibnd), .itxen_in0(vssl_aibnd),
     .itxen_in1(itxen[1]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(odirectin_data_pinp18), .oclkb_in1(vssl_aibnd),
     .odat0_in1(pcs_data_out0_pinp16),
     .odat1_in1(pcs_data_out1_pinp16), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[13]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_pinp18),
     .odat1_aib(odat1_pinp18),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp18),
     .odat0_aib(odat0_pinp18), .oclk_aib(ncdrx_oclk_pinp18),
     .last_bs_out(last_bs_out_pinp18), .oclkb_aib(ncdrx_oclkb_pinp18),
     .jtag_clkdr_in(clkdr_xr7l), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_directout1),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_indat[18]), .oclkn(ncdrx_oclkn_pinp18),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xrx_clkn ( .idata1_in1_jtag_out(idat1_rx_clkn),
     .async_dat_in1_jtag_out(nc_async_dat_rx_clkn),
     .idata0_in1_jtag_out(idat0_rx_clkn),
     .jtag_clkdr_outn(jtag_clkdr_outn_rx_clkn),
     .prev_io_shift_en(rx_shift_en[22]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_rx_clkn),
     .oclk_out(nc_oclk_rx_clkn), .oclkb_out(nc_oclkb_rx_clkn),
     .odat0_out(nc_odat0_out1_rx_clkn),
     .odat1_out(nc_odat1_out1_rx_clkn),
     .odat_async_out(nc_odat_async_out1_rx_clkn),
     .pd_data_out(nc_pd_data_out_rx_clkn), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_l[10]),
     .iclkin_dist_in1(rx_distclk_l[10]), .idata0_in0(vccl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(dft_rx_clk),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .irxen_in1(irxen_r0[2:0]), .istrbclk_in0(rx_strbclk_l[10]),
     .istrbclk_in1(rx_strbclk_l[10]),
     .itxen_in0(idatdll_str_align_stconfig_spare[0]),
     .itxen_in1(vssl_aibnd), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_out0_rx_clkn),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[24]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb),
     .jtag_clkdr_out(nc_jtag_clkdr_out1_rx_clkn),
     .odat1_aib(nc_odat1_out0_rx_clkn),
     .jtag_rx_scan_out(nc_jtag_rx_scan_out1_rx_clkn),
     .odat0_aib(nc_odat0_out0_rx_clkn),
     .oclk_aib(nc_oclk_out0_rx_clkn),
     .last_bs_out(nc_last_bs_out1_rx_clkn),
     .oclkb_aib(nc_oclkb_out0_rx_clkn), .jtag_clkdr_in(clkdr_xr8l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_pinp11),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp11), .iopad(iopad_inclkn),
     .oclkn(oclkn_clkn), .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp11 ( .idata1_in1_jtag_out(nc_idat1_pinp11),
     .async_dat_in1_jtag_out(nc_async_dat_pinp11),
     .idata0_in1_jtag_out(nc_idat0_pinp11),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp11),
     .prev_io_shift_en(rx_shift_en[20]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_pinp11),
     .oclk_out(nc_oclk_pinp11), .oclkb_out(nc_oclkb_pinp11),
     .odat0_out(pcs_data_out0_io[11]),
     .odat1_out(pcs_data_out1_io[11]),
     .odat_async_out(nc_odat_async_pinp11),
     .pd_data_out(nc_pd_data_pinp11), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_l[6]),
     .iclkin_dist_in1(rx_distclk_l[6]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(rx_strbclk_l[6]), .istrbclk_in1(rx_strbclk_l[6]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(nc_odat_async_out0_pinp11),
     .oclkb_in1(vssl_aibnd), .odat0_in1(nc_odat0_out0_rx_clkn),
     .odat1_in1(nc_odat1_out0_rx_clkn), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[22]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_pinp11),
     .odat1_aib(pcs_data_out1_pinp11),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp11),
     .odat0_aib(pcs_data_out0_pinp11), .oclk_aib(nc_oclk_out0_pinp11),
     .last_bs_out(last_bs_out_pinp11),
     .oclkb_aib(nc_oclkb_out0_pinp11), .jtag_clkdr_in(clkdr_xr8l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_pinp13),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp13), .iopad(iopad_indat[11]),
     .oclkn(nc_oclkn_out0_pinp11), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp13 ( .idata1_in1_jtag_out(nc_idat1_pinp13),
     .async_dat_in1_jtag_out(nc_async_dat_pinp13),
     .idata0_in1_jtag_out(nc_idat0_pinp13),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp13),
     .prev_io_shift_en(rx_shift_en[18]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_pinp13),
     .oclk_out(nc_oclk_pinp13), .oclkb_out(nc_oclkb_pinp13),
     .odat0_out(pcs_data_out0_io[13]),
     .odat1_out(pcs_data_out1_io[13]),
     .odat_async_out(nc_odat_async_pinp13),
     .pd_data_out(nc_pd_data_pinp13), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_l[2]),
     .iclkin_dist_in1(rx_distclk_l[2]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(rx_strbclk_l[2]), .istrbclk_in1(rx_strbclk_l[2]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(nc_odat_async_out0_pinp13),
     .oclkb_in1(vssl_aibnd), .odat0_in1(pcs_data_out0_pinp11),
     .odat1_in1(pcs_data_out1_pinp11), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[20]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_pinp13),
     .odat1_aib(pcs_data_out1_pinp13),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp13),
     .odat0_aib(pcs_data_out0_pinp13), .oclk_aib(nc_oclk_out0_pinp13),
     .last_bs_out(last_bs_out_pinp13),
     .oclkb_aib(nc_oclkb_out0_pinp13), .jtag_clkdr_in(clkdr_xr8l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_pinp15),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp15), .iopad(iopad_indat[13]),
     .oclkn(nc_oclkn_out0_pinp13), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp15 ( .idata1_in1_jtag_out(nc_idat1_pinp15),
     .async_dat_in1_jtag_out(nc_async_dat_pinp15),
     .idata0_in1_jtag_out(nc_idat0_pinp15),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp15),
     .prev_io_shift_en(rx_shift_en[16]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_pinp15),
     .oclk_out(nc_oclk_pinp15), .oclkb_out(nc_oclkb_pinp15),
     .odat0_out(pcs_data_out0_io[15]),
     .odat1_out(pcs_data_out1_io[15]),
     .odat_async_out(nc_odat_async_pinp15),
     .pd_data_out(nc_pd_data_pinp15), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_l[0]),
     .iclkin_dist_in1(rx_distclk_l[0]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(rx_strbclk_l[0]), .istrbclk_in1(rx_strbclk_l[0]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(nc_odat_async_out0_pinp15),
     .oclkb_in1(vssl_aibnd), .odat0_in1(pcs_data_out0_pinp13),
     .odat1_in1(pcs_data_out1_pinp13), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[18]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_pinp15),
     .odat1_aib(ncdrx_odat1_pinp15),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp15),
     .odat0_aib(ncdrx_odat0_pinp15), .oclk_aib(ncdrx_oclk_pinp15),
     .last_bs_out(last_bs_out_pinp15), .oclkb_aib(ncdrx_oclkb_pinp15),
     .jtag_clkdr_in(clkdr_xr8l), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_pinp17),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp17), .iopad(iopad_indat[15]),
     .oclkn(ncdrx_oclkn_pinp15), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp17 ( .idata1_in1_jtag_out(nc_idat1_pinp17),
     .async_dat_in1_jtag_out(nc_async_dat_pinp17),
     .idata0_in1_jtag_out(nc_idat0_pinp17),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp17),
     .prev_io_shift_en(rx_shift_en[14]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_pinp17),
     .oclk_out(nc_oclk_pinp17), .oclkb_out(nc_oclkb_pinp17),
     .odat0_out(pcs_data_out0_io[17]),
     .odat1_out(pcs_data_out1_io[17]),
     .odat_async_out(nc_odat_async_pinp17),
     .pd_data_out(nc_pd_data_pinp17), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_l[4]),
     .iclkin_dist_in1(rx_distclk_l[4]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(rx_strbclk_l[4]), .istrbclk_in1(rx_strbclk_l[4]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(nc_odat_async_out0_pinp17),
     .oclkb_in1(vssl_aibnd), .odat0_in1(ncdrx_odat0_pinp15),
     .odat1_in1(ncdrx_odat1_pinp15), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[16]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_pinp17),
     .odat1_aib(pcs_data_out1_pinp17),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp17),
     .odat0_aib(pcs_data_out0_pinp17), .oclk_aib(nc_oclk_out0_pinp17),
     .last_bs_out(last_bs_out_pinp17),
     .oclkb_aib(nc_oclkb_out0_pinp17), .jtag_clkdr_in(clkdr_xr8l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_pinp19),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp19), .iopad(iopad_indat[17]),
     .oclkn(nc_oclkn_out0_pinp17), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp19 ( .idata1_in1_jtag_out(nc_idat1_pinp19),
     .async_dat_in1_jtag_out(nc_async_dat_pinp19),
     .idata0_in1_jtag_out(nc_idat0_pinp19),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp19),
     .prev_io_shift_en(shift_en_outpdir6), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(pd_data_pinp19),
     .oclk_out(nc_oclk_pinp19), .oclkb_out(nc_oclkb_pinp19),
     .odat0_out(pcs_data_out0_io[19]),
     .odat1_out(pcs_data_out1_io[19]),
     .odat_async_out(nc_odat_async_pinp19),
     .pd_data_out(nc_pd_data_pinp19), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(iasync_dat_outpdir6),
     .iclkin_dist_in0(rx_distclk_l[8]), .iclkin_dist_in1(vssl_aibnd),
     .idata0_in0(vssl_aibnd), .idata0_in1(vssl_aibnd),
     .idata1_in0(vssl_aibnd), .idata1_in1(vssl_aibnd),
     .idataselb_in0(vccl_aibnd), .idataselb_in1(idataselb_outpdir6),
     .iddren_in0(vccl_aibnd), .iddren_in1(vssl_aibnd),
     .ilaunch_clk_in0(vssl_aibnd), .ilaunch_clk_in1(vssl_aibnd),
     .ilpbk_dat_in0(vssl_aibnd), .ilpbk_dat_in1(vssl_aibnd),
     .ilpbk_en_in0(vssl_aibnd), .ilpbk_en_in1(vssl_aibnd),
     .indrv_in0({vssl_aibnd, vssl_aibnd}), .indrv_in1(indrv_r78[1:0]),
     .ipdrv_in0({vssl_aibnd, vssl_aibnd}), .ipdrv_in1(ipdrv_r78[1:0]),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .istrbclk_in0(rx_strbclk_l[8]),
     .istrbclk_in1(vssl_aibnd), .itxen_in0(vssl_aibnd),
     .itxen_in1(itxen_outpdir6), .oclk_in1(vssl_aibnd),
     .odat_async_aib(odirectin_data_pinp19), .oclkb_in1(vssl_aibnd),
     .odat0_in1(pcs_data_out0_pinp17),
     .odat1_in1(pcs_data_out1_pinp17), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[14]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_pinp19),
     .odat1_aib(ncdrx_odat1_pinp19),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp19),
     .odat0_aib(ncdrx_odat0_pinp19), .oclk_aib(ncdrx_oclk_pinp19),
     .last_bs_out(last_bs_out_pinp19), .oclkb_aib(ncdrx_oclkb_pinp19),
     .jtag_clkdr_in(clkdr_xr8l), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_outpdir6),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_indat[19]), .oclkn(ncdrx_oclkn_pinp19),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp7 ( .idata1_in1_jtag_out(nc_idat1_pinp7),
     .async_dat_in1_jtag_out(nc_async_dat_pinp7),
     .idata0_in1_jtag_out(nc_idat0_pinp7),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp7),
     .prev_io_shift_en(rx_shift_en[26]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_pinp7),
     .oclk_out(nc_oclk_pinp7), .oclkb_out(nc_oclkb_pinp7),
     .odat0_out(pcs_data_out0_io[7]), .odat1_out(pcs_data_out1_io[7]),
     .odat_async_out(nc_odat_async_pinp7),
     .pd_data_out(nc_pd_data_pinp7), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_r[4]),
     .iclkin_dist_in1(rx_distclk_r[4]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(rx_strbclk_r[4]), .istrbclk_in1(rx_strbclk_r[4]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(nc_odat_async_out0_pinp7),
     .oclkb_in1(vssl_aibnd), .odat0_in1(ncdrx_odat0_pinp5),
     .odat1_in1(ncdrx_odat1_pinp5), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[28]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_pinp7),
     .odat1_aib(pcs_data_out1_pinp7),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp7),
     .odat0_aib(pcs_data_out0_pinp7), .oclk_aib(nc_oclk_out0_pinp7),
     .last_bs_out(last_bs_out_pinp7), .oclkb_aib(nc_oclkb_out0_pinp7),
     .jtag_clkdr_in(clkdr_xr8r), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_pinp9),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp9), .iopad(iopad_indat[7]),
     .oclkn(nc_oclkn_out0_pinp7), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp9 ( .idata1_in1_jtag_out(nc_idat1_pinp9),
     .async_dat_in1_jtag_out(nc_async_dat_pinp9),
     .idata0_in1_jtag_out(nc_idat0_pinp9),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp9),
     .prev_io_shift_en(rx_shift_en[24]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_pinp9),
     .oclk_out(nc_oclk_pinp9), .oclkb_out(nc_oclkb_pinp9),
     .odat0_out(pcs_data_out0_io[9]), .odat1_out(pcs_data_out1_io[9]),
     .odat_async_out(nc_odat_async_pinp9),
     .pd_data_out(nc_pd_data_pinp9), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_r[8]),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(idat0_rx_clkn), .idata1_in0(vssl_aibnd),
     .idata1_in1(idat1_rx_clkn), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vccl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vccl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(dft_rx_clk), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .istrbclk_in0(rx_strbclk_r[8]),
     .istrbclk_in1(vssl_aibnd), .itxen_in0(vssl_aibnd),
     .itxen_in1(vssl_aibnd), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_out0_pinp9), .oclkb_in1(vssl_aibnd),
     .odat0_in1(pcs_data_out0_pinp7), .odat1_in1(pcs_data_out1_pinp7),
     .odat_async_in1(vssl_aibnd), .shift_en(rx_shift_en[26]),
     .pd_data_in1(vssl_aibnd), .dig_rstb(poutp_dig_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_pinp9),
     .odat1_aib(ncdrx_odat1_pinp9),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp9),
     .odat0_aib(ncdrx_odat0_pinp9), .oclk_aib(ncdrx_oclk_pinp9),
     .last_bs_out(last_bs_out_pinp9), .oclkb_aib(ncdrx_oclkb_pinp9),
     .jtag_clkdr_in(clkdr_xr8r), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(nc_jtag_rx_scan_out1_rx_clkn),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(nc_last_bs_out1_rx_clkn), .iopad(iopad_indat[9]),
     .oclkn(oclkn_pinp9), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdirect_in2 (
     .idata1_in1_jtag_out(nc_idat1_directin2),
     .async_dat_in1_jtag_out(nc_async_dat_directin2),
     .idata0_in1_jtag_out(nc_idat0_directin2),
     .jtag_clkdr_outn(jtag_clkdr_outn_directin2),
     .prev_io_shift_en(shift_en_inpshared0),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(input_rstb),
     .pd_data_aib(nc_pd_data_out0_directin[2]),
     .oclk_out(nc_oclk_directin[2]), .oclkb_out(nc_oclkb_directin[2]),
     .odat0_out(nc_odata0_directin[2]),
     .odat1_out(nc_odata1_directin[2]),
     .odat_async_out(odirectin_data[2]),
     .pd_data_out(nc_pd_data_directin[2]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(vssl_aibnd),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vssl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r2[2:0]), .irxen_in1(irxen_inpshared0[2:0]),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odata_async_out0_directin2),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(odat_async_poutp0),
     .shift_en(rx_shift_en[0]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(input_rstb), .jtag_clkdr_out(jtag_clkdr_out_directin2),
     .odat1_aib(nc_odata1_out0_directin[2]),
     .jtag_rx_scan_out(jtag_rx_scan_out_directin2),
     .odat0_aib(nc_odata0_out0_directin[2]), .oclk_aib(oclk_inpdir2),
     .last_bs_out(nc_last_bs_out_directin2), .oclkb_aib(oclkb_inpdir2),
     .jtag_clkdr_in(clkdr_xr3r), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_inpshared0),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_direct_input[2]), .oclkn(nc_oclkn_out0_directin2),
     .iclkn(oclkn_outpdir4_1), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdiin_clkp ( .idata1_in1_jtag_out(nc_idat1_inpclk1),
     .async_dat_in1_jtag_out(nc_async_dat_inpclk1),
     .idata0_in1_jtag_out(nc_idat0_inpclk1),
     .jtag_clkdr_outn(jtag_clkdr_outn_inpclk1),
     .prev_io_shift_en(shift_en_inpdir3), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_diin_clkp),
     .oclk_out(out_rx_fast_clk), .oclkb_out(out_rx_fast_clkb),
     .odat0_out(nc_odat0_diin_clkp), .odat1_out(nc_odat1_diin_clkp),
     .odat_async_out(nc_odat_async_diin_clkp),
     .pd_data_out(nc_pd_data_diin_clkp), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(vssl_aibnd),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vssl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r3[2:0]), .irxen_in1(irxen_inpdir3[2:0]),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(oclk_out0_directin6),
     .odat_async_aib(odat_async_inpclk1),
     .oclkb_in1(oclkb_out0_directin6), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[7]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(input_rstb), .jtag_clkdr_out(jtag_clkdr_out_inpclk1),
     .odat1_aib(nc_odat1_out0_diin_clkp),
     .jtag_rx_scan_out(jtag_rx_scan_out_inpclk1),
     .odat0_aib(nc_odat0_out0_diin_clkp),
     .oclk_aib(nc_oclk_out0_diin_clkp),
     .last_bs_out(nc_last_bs_out_inpclk1),
     .oclkb_aib(nc_oclkb_out0_diin_clkp), .jtag_clkdr_in(clkdr_xr1l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_inpdir3),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_directinclkp), .oclkn(nc_oclkn_out0_diin_clkp),
     .iclkn(rxoclkn_clkn), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdirect_in4 ( .idata1_in1_jtag_out(nc_idat1_inpclk5),
     .async_dat_in1_jtag_out(nc_async_dat_inpclk5),
     .idata0_in1_jtag_out(nc_idat0_inpclk5),
     .jtag_clkdr_outn(jtag_clkdr_outn_inpclk5),
     .prev_io_shift_en(rx_shift_en[1]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_directin[4]),
     .oclk_out(nc_oclk_directin[4]), .oclkb_out(nc_oclkb_directin[4]),
     .odat0_out(nc_odata0_directin[4]),
     .odat1_out(nc_odata1_directin[4]),
     .odat_async_out(odirectin_data[4]),
     .pd_data_out(nc_pd_data_directin[4]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(vssl_aibnd),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vssl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r2[2:0]), .irxen_in1(irxen_r2[2:0]),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(odat_async_inpclk5),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(odat_async_outpclk0),
     .shift_en(rx_shift_en[2]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(input_rstb), .jtag_clkdr_out(jtag_clkdr_out_inpclk5),
     .odat1_aib(nc_odata1_out0_directin[4]),
     .jtag_rx_scan_out(jtag_rx_scan_out_inpclk5),
     .odat0_aib(nc_odata0_out0_directin[4]),
     .oclk_aib(nc_oclk_out0_directin4),
     .last_bs_out(nc_last_bs_out_inptclk5),
     .oclkb_aib(nc_oclkb_out0_directin4), .jtag_clkdr_in(clkdr_xr3l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_inpclk2),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_direct_input[4]), .oclkn(nc_oclkn_out0_directin4),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdout_clkp (
     .idata1_in1_jtag_out(idat1_in0_dout_clkp),
     .async_dat_in1_jtag_out(nc_async_dat_diin_clkp),
     .idata0_in1_jtag_out(idat0_in0_dout_clkp),
     .jtag_clkdr_outn(jtag_clkdr_outn_diin_clkp),
     .prev_io_shift_en(rx_shift_en[2]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_dout_clkp),
     .oclk_out(nc_oclk_dout_clkp), .oclkb_out(nc_oclkb_clkp),
     .odat0_out(nc_odat0_dout_clkp), .odat1_out(nc_odat1_dout_clkp),
     .odat_async_out(nc_odat_async_dout_clkp),
     .pd_data_out(nc_pd_data_dout_clkp), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_diin_clkp),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0_directoutclkp),
     .idata0_in1(vssl_aibnd), .idata1_in0(idat1_directoutclkp),
     .idata1_in1(vssl_aibnd), .idataselb_in0(idataselb[0]),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(txdirclk_fast_clkp),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r34[1:0]),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0(ipdrv_r34[1:0]),
     .ipdrv_in1({vssl_aibnd, vssl_aibnd}), .irxen_in0({vssl_aibnd,
     vccl_aibnd, vssl_aibnd}), .irxen_in1(irxen_r2[2:0]),
     .istrbclk_in0(jtag_clkdr_outn_diin_clkp),
     .istrbclk_in1(vssl_aibnd), .itxen_in0(itxen[0]),
     .itxen_in1(vssl_aibnd), .oclk_in1(oclk_inpclk3),
     .odat_async_aib(odat_async_outpclk0), .oclkb_in1(oclkb_inpclk3),
     .odat0_in1(vssl_aibnd), .odat1_in1(vssl_aibnd),
     .odat_async_in1(vssl_aibnd), .shift_en(rx_shift_en[4]),
     .pd_data_in1(vssl_aibnd), .dig_rstb(input_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_diin_clkp),
     .odat1_aib(nc_odat1_out0_dout_clkp),
     .jtag_rx_scan_out(jtag_rx_scan_out_diin_clkp),
     .odat0_aib(nc_odat0_out0_dout_clkp),
     .oclk_aib(nc_oclk_out0_dout_clkp), .last_bs_out(nc2),
     .oclkb_aib(nc_oclkb_out0_dout_clkp), .jtag_clkdr_in(clkdr_xr3l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_inpclk5),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_directoutclkp), .oclkn(nc_oclkn_out0_dout_clkp),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdirect_in3 ( .idata1_in1_jtag_out(nc_idat1_inpclk6),
     .async_dat_in1_jtag_out(nc_async_dat_inpclk6),
     .idata0_in1_jtag_out(nc_idat0_inpclk6),
     .jtag_clkdr_outn(jtag_clkdr_outn_inpclk6),
     .prev_io_shift_en(shift_en_in_chain1),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(input_rstb),
     .pd_data_aib(nc_pd_data_out0_directin[3]),
     .oclk_out(nc_oclk_directin[3]), .oclkb_out(nc_oclkb_directin[3]),
     .odat0_out(nc_odata0_directin[3]),
     .odat1_out(nc_odata1_directin[3]),
     .odat_async_out(odirectin_data[3]),
     .pd_data_out(nc_pd_data_directin[3]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(vssl_aibnd),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vssl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r2[2:0]), .irxen_in1(irxen_in_chain1[2:0]),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd),
     .odat_async_aib(odirectin_data_out0_chain1),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(odat_async_oshared1),
     .shift_en(rx_shift_en[3]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(input_rstb), .jtag_clkdr_out(jtag_clkdr_inpclk6),
     .odat1_aib(nc_odata1_out0_directin[3]),
     .jtag_rx_scan_out(jtag_rx_scan_inpclk6),
     .odat0_aib(nc_odata0_out0_directin[3]),
     .oclk_aib(nc_oclk_out0_directin3),
     .last_bs_out(last_bs_out_inpclk6),
     .oclkb_aib(nc_oclkb_out0_directin3), .jtag_clkdr_in(clkdr_xr2r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_scan_in_chain1),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_direct_input[3]), .oclkn(nc_oclkn_out0_directin3),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdirect_in5 (
     .idata1_in1_jtag_out(nc_idat1_directin5),
     .async_dat_in1_jtag_out(nc_async_dat_directin5),
     .idata0_in1_jtag_out(nc_idat0_directin5),
     .jtag_clkdr_outn(jtag_clkdr_outn_directin5),
     .prev_io_shift_en(shift_en_inpclk3), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_directin[5]),
     .oclk_out(nc_oclk_directin[5]), .oclkb_out(nc_oclkb_directin[5]),
     .odat0_out(nc_odata0_directin[5]),
     .odat1_out(nc_odata1_directin[5]),
     .odat_async_out(odirectin_data[5]),
     .pd_data_out(nc_pd_data_directin[5]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(vssl_aibnd),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vssl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r2[2:0]), .irxen_in1(irxen_inpclk3[2:0]),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(odat_async_inpclk4),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd),
     .odat_async_in1(nc_odat_async_out0_dout_clkn),
     .shift_en(rx_shift_en[6]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(input_rstb), .jtag_clkdr_out(jtag_clkdr_out_directin5),
     .odat1_aib(nc_odata1_out0_directin[5]),
     .jtag_rx_scan_out(jtag_rx_scan_out_directin5),
     .odat0_aib(nc_odata0_out0_directin[5]),
     .oclk_aib(nc_oclk_out0_directin5),
     .last_bs_out(nc_last_bs_out_outpdir6_1),
     .oclkb_aib(nc_oclkb_out0_directin5), .jtag_clkdr_in(clkdr_xr4l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_inpclk3),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_direct_input[5]), .oclkn(nc_oclkn_inpclk4),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdout_clkn ( .idata1_in1_jtag_out(idat1_dout_clkn),
     .async_dat_in1_jtag_out(nc_async_dat_dout_clkn),
     .idata0_in1_jtag_out(idat0_dout_clkn),
     .jtag_clkdr_outn(jtag_clkdr_outn_dout_clkn),
     .prev_io_shift_en(rx_shift_en[6]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_dout_clkn),
     .oclk_out(nc_oclk_dout_clkn), .oclkb_out(nc_oclkb_clkn),
     .odat0_out(nc_odat0_dout_clkn), .odat1_out(nc_odat1_dout_clkn),
     .odat_async_out(nc_odat_async_dout_clkn),
     .pd_data_out(nc_pd_data_dout_clkn), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_dout_clkn),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0_directoutclkn),
     .idata0_in1(vssl_aibnd), .idata1_in0(idat1_directoutclkn),
     .idata1_in1(vssl_aibnd), .idataselb_in0(idataselb[0]),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(txdirclk_fast_clkn),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r34[1:0]),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0(ipdrv_r34[1:0]),
     .ipdrv_in1({vssl_aibnd, vssl_aibnd}), .irxen_in0({vssl_aibnd,
     vccl_aibnd, vssl_aibnd}), .irxen_in1(irxen_r2[2:0]),
     .istrbclk_in0(jtag_clkdr_outn_dout_clkn),
     .istrbclk_in1(vssl_aibnd), .itxen_in0(itxen[0]),
     .itxen_in1(vssl_aibnd), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_out0_dout_clkn),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[5]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(input_rstb), .jtag_clkdr_out(jtag_clkdr_out_dout_clkn),
     .odat1_aib(nc_odat1_out0_dout_clkn),
     .jtag_rx_scan_out(jtag_rx_scan_out_dout_clkn),
     .odat0_aib(nc_odat0_out0_dout_clkn),
     .oclk_aib(nc_oclk_out0_dout_clkn),
     .last_bs_out(nc_last_bs_out_dout_clkn),
     .oclkb_aib(nc_oclkb_out0_dout_clkn), .jtag_clkdr_in(clkdr_xr4l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_directin5),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_directoutclkn), .oclkn(nc_oclkn_out0_dout_clkn),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdirect_out0 (
     .idata1_in1_jtag_out(nc_idat1_outpclk1_1),
     .async_dat_in1_jtag_out(async_dat_outpclk1_1),
     .idata0_in1_jtag_out(nc_idat0_outpclk1_1),
     .jtag_clkdr_outn(jtag_clkdr_outn_outpclk1_1),
     .prev_io_shift_en(shift_en_vinp0), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb),
     .pd_data_aib(nc_pd_data_out0_directout[0]),
     .oclk_out(nc_oclk_directout[0]),
     .oclkb_out(nc_oclkb_directout[0]),
     .odat0_out(nc_odat0_directout[0]),
     .odat1_out(nc_odat1_directout[0]),
     .odat_async_out(nc_odat_async_directout[0]),
     .pd_data_out(nc_pd_data_directout[0]),
     .async_dat_in0(idirectout_data[0]), .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(iclkin_dist_vinp0),
     .iclkin_dist_in1(iclkin_dist_vinp0), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(idataselb[1]),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r12[1:0]),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0(ipdrv_r12[1:0]),
     .ipdrv_in1({vssl_aibnd, vssl_aibnd}), .irxen_in0({vssl_aibnd,
     vccl_aibnd, vssl_aibnd}), .irxen_in1(irxen_vinp0[2:0]),
     .istrbclk_in0(istrbclk_vinp0), .istrbclk_in1(istrbclk_vinp0),
     .itxen_in0(itxen[1]), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_out0_directout[0]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[10]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(avmm_sync_rstb), .jtag_clkdr_out(jtag_clkdr_outpclk1_1),
     .odat1_aib(odat1_outpclk1_1),
     .jtag_rx_scan_out(jtag_rx_scan_outpclk1_1),
     .odat0_aib(odat0_outpclk1_1),
     .oclk_aib(nc_oclk_out0_directout[0]),
     .last_bs_out(nc_last_bs_out_directout0),
     .oclkb_aib(nc_oclkb_out0_directout[0]),
     .jtag_clkdr_in(clkdr_xr1l), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_vinp0),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_directout[0]), .oclkn(nc_oclkn_out0_directout[0]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp5 ( .idata1_in1_jtag_out(nc_idat1_pinp5),
     .async_dat_in1_jtag_out(nc_async_dat_pinp5),
     .idata0_in1_jtag_out(nc_idat0_pinp5),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp5),
     .prev_io_shift_en(rx_shift_en[28]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_pinp5),
     .oclk_out(nc_oclk_pinp5), .oclkb_out(nc_oclkb_pinp5),
     .odat0_out(pcs_data_out0_io[5]), .odat1_out(pcs_data_out1_io[5]),
     .odat_async_out(nc_odat_async_pinp5),
     .pd_data_out(nc_pd_data_pinp5), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_r[0]),
     .iclkin_dist_in1(rx_distclk_r[0]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(rx_strbclk_r[0]), .istrbclk_in1(rx_strbclk_r[0]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(nc_odat_async_out0_pinp5),
     .oclkb_in1(vssl_aibnd), .odat0_in1(pcs_data_out0_pinp3),
     .odat1_in1(pcs_data_out1_pinp3), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[30]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_pinp5),
     .odat1_aib(ncdrx_odat1_pinp5),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp5),
     .odat0_aib(ncdrx_odat0_pinp5), .oclk_aib(ncdrx_oclk_pinp5),
     .last_bs_out(last_bs_out_pinp5), .oclkb_aib(ncdrx_oclkb_pinp5),
     .jtag_clkdr_in(clkdr_xr8r), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_pinp7),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp7), .test_weakpd(jtag_weakpdn),
     .test_weakpu(jtag_weakpu), .iopad(iopad_indat[5]),
     .oclkn(ncdrx_oclkn_pinp5), .iclkn(vssl_aibnd));
aibnd_buffx1_top xdirect_out2 ( .idata1_in1_jtag_out(nc_idat1_dirout2),
     .async_dat_in1_jtag_out(idirectout_data_outpdir2_1),
     .idata0_in1_jtag_out(nc_idat0_dirout2),
     .jtag_clkdr_outn(jtag_clkdr_outn_dirout2),
     .prev_io_shift_en(rx_shift_en[5]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb),
     .pd_data_aib(nc_pd_data_out0_directout[2]),
     .oclk_out(nc_oclk_directout[2]),
     .oclkb_out(nc_oclkb_directout[2]),
     .odat0_out(nc_odat0_directout[2]),
     .odat1_out(nc_odat1_directout[2]),
     .odat_async_out(nc_odat_async_directout[2]),
     .pd_data_out(nc_pd_data_directout[2]),
     .async_dat_in0(idirectout_data[2]), .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(vssl_aibnd), .iclkin_dist_in1(vssl_aibnd),
     .idata0_in0(vssl_aibnd), .idata0_in1(idat0_dout_clkn),
     .idata1_in0(vssl_aibnd), .idata1_in1(idat1_dout_clkn),
     .idataselb_in0(idataselb[1]), .idataselb_in1(idataselb[0]),
     .iddren_in0(vssl_aibnd), .iddren_in1(vccl_aibnd),
     .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(txdirclk_fast_clkn), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r34[1:0]),
     .indrv_in1(indrv_r34[1:0]), .ipdrv_in0(ipdrv_r34[1:0]),
     .ipdrv_in1(ipdrv_r34[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(vssl_aibnd), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[1]), .itxen_in1(itxen[0]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_out0_directout[2]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[9]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(input_rstb), .jtag_clkdr_out(jtag_clkdr_out_dirout2),
     .odat1_aib(nc_odat1_out0_directout[2]),
     .jtag_rx_scan_out(jtag_rx_scan_out_dirout2),
     .odat0_aib(nc_odat0_out0_directout[2]),
     .oclk_aib(nc_oclk_out0_directout[2]),
     .last_bs_out(nc_last_bs_out_dirout2),
     .oclkb_aib(nc_oclkb_out0_directout[2]),
     .jtag_clkdr_in(clkdr_xr4l), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_dout_clkn),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_directout[2]), .oclkn(nc_oclkn_out0_directout[2]),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdiin_clkn ( .idata1_in1_jtag_out(nc_idat1_inpclk1n),
     .async_dat_in1_jtag_out(nc_async_dat_inpclk1n),
     .idata0_in1_jtag_out(nc_idat0_inpclk1n),
     .jtag_clkdr_outn(jtag_clkdr_outn_inpclk1n),
     .prev_io_shift_en(rx_shift_en[35]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_diin_clkn),
     .oclk_out(nc_oclk_diin_clkn), .oclkb_out(nc_oclkb_diin_clkn),
     .odat0_out(nc_odat0_diin_clkn), .odat1_out(nc_odat1_diin_clkn),
     .odat_async_out(nc_odat_async_diin_clkn),
     .pd_data_out(nc_pd_data_diin_clkn), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(vssl_aibnd),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vssl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .irxen_in1(irxen_r2[2:0]), .istrbclk_in0(vssl_aibnd),
     .istrbclk_in1(vssl_aibnd), .itxen_in0(vssl_aibnd),
     .itxen_in1(vssl_aibnd), .oclk_in1(vssl_aibnd),
     .odat_async_aib(odat_async_out_inpclk1n), .oclkb_in1(vssl_aibnd),
     .odat0_in1(vssl_aibnd), .odat1_in1(vssl_aibnd),
     .odat_async_in1(vssl_aibnd), .shift_en(rx_shift_en[8]),
     .pd_data_in1(vssl_aibnd), .dig_rstb(input_rstb),
     .jtag_clkdr_out(jtag_clkdr_inpclk1n),
     .odat1_aib(nc_odat1_out0_diin_clkn),
     .jtag_rx_scan_out(jtag_rx_scan_inpclk1n),
     .odat0_aib(nc_odat0_out0_diin_clkn),
     .oclk_aib(nc_oclk_out0_diin_clkn),
     .last_bs_out(last_bs_out_inpclk1n),
     .oclkb_aib(nc_oclkb_out0_diin_clkn), .jtag_clkdr_in(clkdr_xr2l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_inpdir4),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_directinclkn), .oclkn(rxoclkn_clkn),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp3 ( .idata1_in1_jtag_out(nc_idat1_pinp3),
     .async_dat_in1_jtag_out(nc_async_dat_pinp3),
     .idata0_in1_jtag_out(nc_idat0_pinp3),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp3),
     .prev_io_shift_en(rx_shift_en[30]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_pinp3),
     .oclk_out(nc_oclk_pinp3), .oclkb_out(nc_oclkb_pinp3),
     .odat0_out(pcs_data_out0_io[3]), .odat1_out(pcs_data_out1_io[3]),
     .odat_async_out(nc_odat_async_pinp3),
     .pd_data_out(nc_pd_data_pinp3), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_r[2]),
     .iclkin_dist_in1(rx_distclk_r[2]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(rx_strbclk_r[2]), .istrbclk_in1(rx_strbclk_r[2]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(nc_odat_async_out0_pinp3),
     .oclkb_in1(vssl_aibnd), .odat0_in1(pcs_data_out0_pinp1),
     .odat1_in1(pcs_data_out1_pinp1), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[32]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_pinp3),
     .odat1_aib(pcs_data_out1_pinp3),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp3),
     .odat0_aib(pcs_data_out0_pinp3), .oclk_aib(nc_oclk_out0_pinp3),
     .last_bs_out(last_bs_out_pinp3), .oclkb_aib(nc_oclkb_out0_pinp3),
     .jtag_clkdr_in(clkdr_xr8r), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_pinp5),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp5), .iopad(iopad_indat[3]),
     .oclkn(nc_oclkn_out0_pinp3), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xpinp1 ( .idata1_in1_jtag_out(nc_idat1_pinp1),
     .async_dat_in1_jtag_out(nc_async_dat_pinp1),
     .idata0_in1_jtag_out(nc_idat0_pinp1),
     .jtag_clkdr_outn(jtag_clkdr_outn_pinp1),
     .prev_io_shift_en(rx_shift_en[32]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_pinp1),
     .oclk_out(nc_oclk_pinp1), .oclkb_out(nc_oclkb_pinp1),
     .odat0_out(pcs_data_out0_io[1]), .odat1_out(pcs_data_out1_io[1]),
     .odat_async_out(nc_odat_async_pinp1),
     .pd_data_out(nc_pd_data_pinp1), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_r[6]),
     .iclkin_dist_in1(rx_distclk_r[6]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r0[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(rx_strbclk_r[6]), .istrbclk_in1(rx_strbclk_r[6]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(nc_odat_async_out0_pinp1),
     .oclkb_in1(vssl_aibnd), .odat0_in1(nc_odata0_out0_directin[1]),
     .odat1_in1(nc_odata1_out0_directin[1]),
     .odat_async_in1(vssl_aibnd), .shift_en(rx_shift_en[34]),
     .pd_data_in1(vssl_aibnd), .dig_rstb(poutp_dig_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_pinp1),
     .odat1_aib(pcs_data_out1_pinp1),
     .jtag_rx_scan_out(jtag_rx_scan_out_pinp1),
     .odat0_aib(pcs_data_out0_pinp1), .oclk_aib(nc_oclk_out0_pinp1),
     .last_bs_out(last_bs_out_pinp1), .oclkb_aib(nc_oclkb_out0_pinp1),
     .jtag_clkdr_in(clkdr_xr8r), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_pinp3),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp3), .test_weakpd(jtag_weakpdn),
     .test_weakpu(jtag_weakpu), .iopad(iopad_indat[1]),
     .oclkn(nc_oclkn_out0_pinp1), .iclkn(vssl_aibnd));
aibnd_buffx1_top xdirect_in0 ( .idata1_in1_jtag_out(nc_idat1_inpdir4),
     .async_dat_in1_jtag_out(nc_async_dat_inpdir4),
     .idata0_in1_jtag_out(nc_idat0_inpdir4),
     .jtag_clkdr_outn(jtag_clkdr_outn_inpdir4),
     .prev_io_shift_en(shift_en_inpclk0n), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_directin[0]),
     .oclk_out(nc_oclk_directin[0]), .oclkb_out(nc_oclkb_directin[0]),
     .odat0_out(nc_odata0_directin[0]),
     .odat1_out(nc_odata1_directin[0]),
     .odat_async_out(odirectin_data[0]),
     .pd_data_out(nc_pd_data_directin[0]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(vssl_aibnd),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vssl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r2[2:0]), .irxen_in1({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .istrbclk_in0(vssl_aibnd),
     .istrbclk_in1(vssl_aibnd), .itxen_in0(vssl_aibnd),
     .itxen_in1(vssl_aibnd), .oclk_in1(vssl_aibnd),
     .odat_async_aib(odirectin_data_out0[0]), .oclkb_in1(vssl_aibnd),
     .odat0_in1(vssl_aibnd), .odat1_in1(vssl_aibnd),
     .odat_async_in1(odat_async_out_inpclk1n),
     .shift_en(rx_shift_en[35]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb),
     .jtag_clkdr_out(jtag_clkdr_out_inpdir4),
     .odat1_aib(nc_odat1_directin0),
     .jtag_rx_scan_out(jtag_rx_scan_out_inpdir4),
     .odat0_aib(nc_odat0_directin0),
     .oclk_aib(nc_oclk_out0_directin[0]),
     .last_bs_out(last_bs_out_inpdir4),
     .oclkb_aib(nc_oclkb_out0_directin[0]), .jtag_clkdr_in(clkdr_xr2l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_inpclk0n),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_direct_input[0]), .oclkn(oclkn_inpdir4),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xdirect_in1 ( .idata1_in1_jtag_out(nc_idat1_inpdir1),
     .async_dat_in1_jtag_out(nc_async_dat_inpdir1),
     .idata0_in1_jtag_out(nc_idat0_inpdir1),
     .jtag_clkdr_outn(jtag_clkdr_outn_inpdir1),
     .prev_io_shift_en(rx_shift_en[34]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(input_rstb), .pd_data_aib(nc_pd_data_out0_directin[1]),
     .oclk_out(nc_oclk_directin[1]), .oclkb_out(nc_oclkb_directin[1]),
     .odat0_out(nc_odata0_directin[1]),
     .odat1_out(nc_odata1_directin[1]),
     .odat_async_out(odirectin_data[1]),
     .pd_data_out(nc_pd_data_directin[1]), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_r[10]),
     .iclkin_dist_in1(rx_distclk_r[10]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vssl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r2[2:0]), .irxen_in1(irxen_r0[2:0]),
     .istrbclk_in0(rx_strbclk_r[10]), .istrbclk_in1(rx_strbclk_r[10]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(odirectin_data_out0[1]),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(odirectin_data_in_chain1),
     .shift_en(rx_shift_en[36]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(poutp_dig_rstb), .jtag_clkdr_out(jtag_clkdr_out_chain1),
     .odat1_aib(nc_odata1_out0_directin[1]),
     .jtag_rx_scan_out(jtag_scan_out_chain1),
     .odat0_aib(nc_odata0_out0_directin[1]),
     .oclk_aib(nc_oclk_out0_directin[1]),
     .last_bs_out(last_bs_out_chain1),
     .oclkb_aib(nc_oclkb_out0_directin[1]), .jtag_clkdr_in(clkdr_xr8r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_pinp1),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_pinp1), .iopad(iopad_direct_input[1]),
     .oclkn(nc_oclkn_out0_directin[1]), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_str_align x982 ( .vcc_aibnd(vccl_aibnd), .vss_aibnd(vssl_aibnd),
     .scan_shift_n(idatdll_scan_shift_n),
     .rb_clkdiv_str(idatdll_rb_clkdiv_str[2:0]),
     .scan_rst_n(idatdll_scan_rst_n), .ref_clk_p(oclk_clkp),
     .lstrbclk_l_11(rx_strbclk_l[11]), .vcc_io(vccl_aibnd),
     .lstrbclk_l_10(rx_strbclk_l[10]),
     .odll_dll2core_str(odll_dll2core_str[12:0]),
     .lstrbclk_l_9(rx_strbclk_l[9]), .lstrbclk_l_8(rx_strbclk_l[8]),
     .lstrbclk_l_7(rx_strbclk_l[7]), .lstrbclk_l_6(rx_strbclk_l[6]),
     .lstrbclk_l_5(rx_strbclk_l[5]), .lstrbclk_l_4(rx_strbclk_l[4]),
     .lstrbclk_l_3(rx_strbclk_l[3]), .lstrbclk_l_2(rx_strbclk_l[2]),
     .lstrbclk_l_1(rx_strbclk_l[1]), .lstrbclk_l_0(rx_strbclk_l[0]),
     .lstrbclk_r_0(rx_strbclk_r[0]), .lstrbclk_r_1(rx_strbclk_r[1]),
     .lstrbclk_r_2(rx_strbclk_r[2]),
     .idll_core2dll_str(idll_core2dll_str[2:0]),
     .lstrbclk_r_3(rx_strbclk_r[3]), .idll_lock_req(idll_lock_req),
     .idll_entest_str(idatdll_entest_str),
     .lstrbclk_r_4(rx_strbclk_r[4]), .lstrbclk_r_5(rx_strbclk_r[5]),
     .lstrbclk_r_6(rx_strbclk_r[6]), .lstrbclk_r_7(rx_strbclk_r[7]),
     .lstrbclk_r_8(rx_strbclk_r[8]), .lstrbclk_r_9(rx_strbclk_r[9]),
     .lstrbclk_r_10(rx_strbclk_r[10]),
     .lstrbclk_r_11(rx_strbclk_r[11]),
     .scan_mode_n(idatdll_scan_mode_n),
     .pipeline_global_en(idatdll_pipeline_global_en),
     .scan_clk_in(idatdll_scan_clk_in), .scan_in(idatdll_scan_in),
     .scan_out(dll_scan_out), .csr_reg_str(csr_reg_str[51:0]),
     .odll_lock(odll_lock),
     .rb_half_code_str(idatdll_rb_half_code_str),
     .rb_selflock_str(idatdll_rb_selflock_str), .ref_clk_n(oclk_clkpb),
     .test_clk_pll_en_n(idatdll_test_clk_pll_en_n));

aibnd_clkmux2 xrx_clkp_mux ( 
      .oclk_out(oclk_clkp),
     .mux_sel(rx_shift_en[23]), .oclk_in0(drx_oclk_out0_rx_clkp),
     .oclk_in1(oclk_pinp8));

aibnd_clkmux2 xrx_clkn_mux ( 
      .oclk_out(oclk_clkpb),
     .mux_sel(rx_shift_en[23]), .oclk_in0(drx_oclkb_out0_rx_clkp),
     .oclk_in1(oclkb_pinp8));

assign oclk_clkp_buf = oclk_clkp;
assign oclk_clkpb_buf = oclk_clkpb;

assign scan_out = dll_scan_out;
assign pcs_data_out0[3] = pcs_data_out0_io[3];
assign pcs_data_out0[5] = pcs_data_out0_io[5];
assign pcs_data_out1[5] = pcs_data_out1_io[5];
assign pcs_data_out1[7] = pcs_data_out1_io[7];
assign pcs_data_out0[7] = pcs_data_out0_io[7];
assign pcs_data_out0[9] = pcs_data_out0_io[9];
assign pcs_data_out1[9] = pcs_data_out1_io[9];
assign pcs_data_out0[11] = pcs_data_out0_io[11];
assign pcs_data_out1[11] = pcs_data_out1_io[11];
assign pcs_data_out1[13] = pcs_data_out1_io[13];
assign pcs_data_out0[13] = pcs_data_out0_io[13];
assign pcs_data_out0[15] = pcs_data_out0_io[15];
assign pcs_data_out1[15] = pcs_data_out1_io[15];
assign pcs_data_out1[17] = pcs_data_out1_io[17];
assign pcs_data_out0[17] = pcs_data_out0_io[17];
assign pcs_data_out0[19] = pcs_data_out0_io[19];
assign pcs_data_out1[19] = pcs_data_out1_io[19];
assign pcs_data_out0[0] = pcs_data_out0_io[0];
assign pcs_data_out1[0] = pcs_data_out1_io[0];
assign pcs_data_out1[2] = pcs_data_out1_io[2];
assign pcs_data_out0[2] = pcs_data_out0_io[2];
assign pcs_data_out0[4] = pcs_data_out0_io[4];
assign pcs_data_out1[4] = pcs_data_out1_io[4];
assign pcs_data_out1[6] = pcs_data_out1_io[6];
assign pcs_data_out0[6] = pcs_data_out0_io[6];
assign pcs_data_out0[8] = pcs_data_out0_io[8];
assign pcs_data_out1[8] = pcs_data_out1_io[8];
assign pcs_data_out1[10] = pcs_data_out1_io[10];
assign pcs_data_out0[10] = pcs_data_out0_io[10];
assign pcs_data_out0[12] = pcs_data_out0_io[12];
assign pcs_data_out1[12] = pcs_data_out1_io[12];
assign pcs_data_out1[14] = pcs_data_out1_io[14];
assign pcs_data_out0[14] = pcs_data_out0_io[14];
assign pcs_data_out0[16] = pcs_data_out0_io[16];
assign pcs_data_out1[16] = pcs_data_out1_io[16];
assign pcs_data_out0[18] = pcs_data_out0_io[18];
assign pcs_data_out1[18] = pcs_data_out1_io[18];
assign pcs_data_out0[1] = pcs_data_out0_io[1];
assign pcs_data_out1[3] = pcs_data_out1_io[3];
assign pcs_data_out1[1] = pcs_data_out1_io[1];

assign pre_pcs_clk = pcs_clk_inv;

assign pcs_clk_inv = lstrbclk_rep;
aibnd_rxdat_mimic x1231 ( .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .odat_out(pcs_clk),
     .odat_in(pre_pcs_clk));

endmodule

