// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. All rights reserved
`ifndef c3dfx_dv_vh
`define c3dfx_dv_vh

`define C3DFX_RTL_MODE

`endif // c3dfx_dv_vh

