// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. All rights reserved
wire [79:0] pld_rx_fabric_data_out;
ndaibadapt_wrap  ndut(

// EMIB inout
                      .io_aib0(aib0), 
                      .io_aib1(aib1), 
                      .io_aib10(aib10),
                      .io_aib11(aib11),
                      .io_aib12(aib12),
                      .io_aib13(aib13),
                      .io_aib14(aib14),
                      .io_aib15(aib15),
                      .io_aib16(aib16),
                      .io_aib17(aib17),
                      .io_aib18(aib18),
                      .io_aib19(aib19),
                      .io_aib2(aib2), 
                      .io_aib20(aib20),
                      .io_aib21(aib21),
                      .io_aib22(aib22),
                      .io_aib23(aib23),
                      .io_aib24(aib24),
                      .io_aib25(aib25),
                      .io_aib26(aib26),
                      .io_aib27(aib27),
                      .io_aib28(aib28),
                      .io_aib29(aib29),
                      .io_aib3(aib3), 
                      .io_aib30(aib30),
                      .io_aib31(aib31),
                      .io_aib32(aib32),
                      .io_aib33(aib33),
                      .io_aib34(aib34),
                      .io_aib35(aib35),
                      .io_aib36(aib36),
                      .io_aib37(aib37),
                      .io_aib38(aib38),
                      .io_aib39(aib39),
                      .io_aib4(aib4), 
                      .io_aib40(aib40),
                      .io_aib41(aib41),
                      .io_aib42(aib42),
                      .io_aib43(aib43),
                      .io_aib44(aib44),
                      .io_aib45(aib45),
                      .io_aib46(aib46),
                      .io_aib47(aib47),
                      .io_aib48(aib48),
                      .io_aib49(aib49),
                      .io_aib5(aib5), 
                      .io_aib50(aib50),
                      .io_aib51(aib51),
                      .io_aib52(aib52),
                      .io_aib53(aib53),
                      .io_aib54(aib54),
                      .io_aib55(aib55),
                      .io_aib56(aib56),
                      .io_aib57(aib57),
                      .io_aib58(aib58),
                      .io_aib59(aib59),
                      .io_aib6(aib6), 
                      .io_aib60(aib60),
                      .io_aib61(aib61),
                      .io_aib62(aib62),
                      .io_aib63(aib63),
                      .io_aib64(aib64),
                      .io_aib65(aib65),
                      .io_aib66(aib66),
                      .io_aib67(aib67),
                      .io_aib68(aib68),
                      .io_aib69(aib69),
                      .io_aib7(aib7), 
                      .io_aib70(aib70),
                      .io_aib71(aib71),
                      .io_aib72(aib72),
                      .io_aib73(aib73),
                      .io_aib74(aib74),
                      .io_aib75(aib75),
                      .io_aib76(aib76),
                      .io_aib77(aib77),
                      .io_aib78(aib78),
                      .io_aib79(aib79),
                      .io_aib8(aib8), 
                      .io_aib80(aib80),
                      .io_aib81(aib81),
                      .io_aib82(aib82),
                      .io_aib83(aib83),
                      .io_aib84(aib84),
                      .io_aib85(aib85),
                      .io_aib86(aib86),
                      .io_aib87(aib87),
                      .io_aib88(aib88),
                      .io_aib89(aib89),
                      .io_aib9(aib9), 
                      .io_aib90(aib90),
                      .io_aib91(aib91),
                      .io_aib92(aib92),
                      .io_aib93(aib93),
                      .io_aib94(aib94),
                      .io_aib95(aib95),

    // Adapter       input 
              	      .bond_rx_asn_ds_in_fifo_hold(1'b0),
              	      .bond_rx_asn_us_in_fifo_hold(1'b0),
              	      .bond_rx_fifo_ds_in_rden(1'b0),
              	      .bond_rx_fifo_ds_in_wren(1'b0),
              	      .bond_rx_fifo_us_in_rden(1'b0),
              	      .bond_rx_fifo_us_in_wren(1'b0),
                      .bond_rx_hrdrst_ds_in_fabric_rx_dll_lock(1'b0),
                      .bond_rx_hrdrst_us_in_fabric_rx_dll_lock(1'b0),
                      .bond_rx_hrdrst_ds_in_fabric_rx_dll_lock_req(1'b0),
                      .bond_rx_hrdrst_us_in_fabric_rx_dll_lock_req(1'b0),
              	      .bond_tx_fifo_ds_in_dv(1'b0),
              	      .bond_tx_fifo_ds_in_rden(1'b0),
              	      .bond_tx_fifo_ds_in_wren(1'b0),
              	      .bond_tx_fifo_us_in_dv(1'b0),
              	      .bond_tx_fifo_us_in_rden(1'b0),
              	      .bond_tx_fifo_us_in_wren(1'b0),
                      .bond_tx_hrdrst_ds_in_fabric_tx_dcd_cal_done(1'b0),
                      .bond_tx_hrdrst_us_in_fabric_tx_dcd_cal_done(1'b0),
                      .bond_tx_hrdrst_ds_in_fabric_tx_dcd_cal_req(1'b0),
                      .bond_tx_hrdrst_us_in_fabric_tx_dcd_cal_req(1'b0),
    
    // Config  input 
                      .csr_config(csr_config),
                      .csr_clk_in(csr_clk_in),
                      .csr_in(csr_in),
                      .csr_pipe_in(csr_pipe_in),
                      .csr_rdy_dly_in(csr_rdy_dly_in),
                      .csr_rdy_in(csr_rdy_in),
                      .nfrzdrv_in(nfrzdrv_in),
                      .usermode_in(usermode_in),
    
    // PLD input
              	      .hip_aib_fsr_in(hip_aib_fsr_in),
              	      .hip_aib_ssr_in(hip_aib_ssr_in),
              	      .hip_avmm_read(hip_avmm_read),
              	      .hip_avmm_reg_addr(hip_avmm_reg_addr),
              	      .hip_avmm_write(hip_avmm_write),
              	      .hip_avmm_writedata(hip_avmm_writedata),
              	      .pld_10g_krfec_rx_clr_errblk_cnt(pld_10g_krfec_rx_clr_errblk_cnt),
              	      .pld_10g_rx_align_clr(pld_10g_rx_align_clr),
              	      .pld_10g_rx_clr_ber_count(pld_10g_rx_clr_ber_count),
              	      .pld_10g_tx_bitslip(pld_10g_tx_bitslip),
              	      .pld_10g_tx_burst_en(pld_10g_tx_burst_en),
              	      .pld_10g_tx_diag_status(pld_10g_tx_diag_status),
              	      .pld_10g_tx_wordslip(pld_10g_tx_wordslip),
              	      .pld_8g_a1a2_size(pld_8g_a1a2_size),
              	      .pld_8g_bitloc_rev_en(pld_8g_bitloc_rev_en),
              	      .pld_8g_byte_rev_en(pld_8g_byte_rev_en),
              	      .pld_8g_eidleinfersel(pld_8g_eidleinfersel),
              	      .pld_8g_encdt(pld_8g_encdt),
              	      .pld_8g_tx_boundary_sel(pld_8g_tx_boundary_sel),
              	      .pld_adapter_rx_pld_rst_n(pld_adapter_rx_pld_rst_n),
              	      .pld_adapter_tx_pld_rst_n(pld_adapter_tx_pld_rst_n),
              	      .pld_avmm1_clk_rowclk(pld_avmm1_clk_rowclk),
              	      .pld_avmm1_read(pld_avmm1_read),
              	      .pld_avmm1_reg_addr(pld_avmm1_reg_addr),
              	      .pld_avmm1_request(pld_avmm1_request),
              	      .pld_avmm1_write(pld_avmm1_write),
              	      .pld_avmm1_writedata(pld_avmm1_writedata),
              	      .pld_avmm1_reserved_in(pld_avmm1_reserved_in),
              	      .pld_avmm2_clk_rowclk(pld_avmm2_clk_rowclk),
              	      .pld_avmm2_read(pld_avmm2_read),
              	      .pld_avmm2_reg_addr(pld_avmm2_reg_addr),
              	      .pld_avmm2_request(pld_avmm2_request),
              	      .pld_avmm2_write(pld_avmm2_write),
              	      .pld_avmm2_writedata(pld_avmm2_writedata),
              	      .pld_avmm2_reserved_in(pld_avmm2_reserved_in),
              	      .pld_bitslip(pld_bitslip),
              	      .pld_fpll_shared_direct_async_in(pld_fpll_shared_direct_async_in),
              	      .pld_fpll_shared_direct_async_in_rowclk(pld_fpll_shared_direct_async_in_rowclk),
              	      .pld_fpll_shared_direct_async_in_dcm(pld_fpll_shared_direct_async_in_dcm),
              	      .pld_ltr(pld_ltr),
              	      .pr_channel_freeze_n(pr_channel_freeze_n),
              	      .pld_pcs_rx_pld_rst_n(pld_pcs_rx_pld_rst_n),
              	      .pld_pcs_tx_pld_rst_n(pld_pcs_tx_pld_rst_n),
              	      .pld_pma_adapt_start(pld_pma_adapt_start),
              	      .pld_pma_coreclkin_rowclk(pld_pma_coreclkin_rowclk),
              	      .pld_pma_csr_test_dis(pld_pma_csr_test_dis),
              	      .pld_pma_early_eios(pld_pma_early_eios),
              	      .pld_pma_eye_monitor(pld_pma_eye_monitor),
              	      .pld_pma_fpll_cnt_sel(pld_pma_fpll_cnt_sel),
              	      .pld_pma_fpll_extswitch(pld_pma_fpll_extswitch),
              	      .pld_pma_fpll_lc_csr_test_dis(pld_pma_fpll_lc_csr_test_dis),
              	      .pld_pma_fpll_num_phase_shifts(pld_pma_fpll_num_phase_shifts),
              	      .pld_pma_fpll_pfden(pld_pma_fpll_pfden),
              	      .pld_pma_fpll_up_dn_lc_lf_rstn(pld_pma_fpll_up_dn_lc_lf_rstn),
              	      .pld_pma_ltd_b(pld_pma_ltd_b),
              	      .pld_pma_nrpi_freeze(pld_pma_nrpi_freeze),
              	      .pld_pma_pcie_switch(pld_pma_pcie_switch),
              	      .pld_pma_ppm_lock(pld_pma_ppm_lock),
              	      .pld_pma_reserved_out(pld_pma_reserved_out),
              	      .pld_pma_rs_lpbk_b(pld_pma_rs_lpbk_b),
              	      .pld_pma_rxpma_rstb(pld_pma_rxpma_rstb),
              	      .pld_pma_tx_bitslip(pld_pma_tx_bitslip),
              	      .pld_pma_txdetectrx(pld_pma_txdetectrx),
              	      .pld_pma_txpma_rstb(pld_pma_txpma_rstb),
              	      .pld_pmaif_rxclkslip(pld_pmaif_rxclkslip),
              	      .pld_polinv_rx(pld_polinv_rx),
              	      .pld_polinv_tx(pld_polinv_tx),
              	      .pld_rx_clk1_rowclk(pld_rx_clk1_rowclk),
              	      .pld_rx_clk2_rowclk(pld_rx_clk2_rowclk),
              	      .pld_rx_dll_lock_req(pld_rx_dll_lock_req),
              	      .pld_rx_fabric_fifo_align_clr(pld_rx_fabric_fifo_align_clr),
              	      .pld_rx_fabric_fifo_rd_en(pld_rx_fabric_fifo_rd_en),
              	      .pld_rx_prbs_err_clr(pld_rx_prbs_err_clr),
              	      .pld_sclk1_rowclk(pld_sclk1_rowclk),
              	      .pld_sclk2_rowclk(pld_sclk2_rowclk),
              	      .pld_syncsm_en(pld_syncsm_en),
              	      .pld_tx_clk1_rowclk(pld_rx_clk1_rowclk),
              	      .pld_tx_clk2_rowclk(pld_rx_clk2_rowclk),
              	      .pld_tx_fabric_data_in(pld_rx_fabric_data_out),  //Loopback from rx
              	      .pld_txelecidle(pld_txelecidle),
                      .pld_tx_dll_lock_req(pld_tx_dll_lock_req),
                      .pld_tx_fifo_latency_adj_en(pld_tx_fifo_latency_adj_en),
                      .pld_rx_fifo_latency_adj_en(pld_rx_fifo_latency_adj_en),
                      .pld_aib_fabric_rx_dll_lock_req(pld_aib_fabric_rx_dll_lock_req),
                      .pld_aib_fabric_tx_dcd_cal_req(pld_aib_fabric_tx_dcd_cal_req),
                      .pld_aib_hssi_tx_dcd_cal_req(pld_aib_hssi_tx_dcd_cal_req),
                      .pld_aib_hssi_tx_dll_lock_req(pld_aib_hssi_tx_dll_lock_req),
                      .pld_aib_hssi_rx_dcd_cal_req(pld_aib_hssi_rx_dcd_cal_req),
                      .pld_tx_ssr_reserved_in(pld_tx_ssr_reserved_in), 
                      .pld_rx_ssr_reserved_in(pld_rx_ssr_reserved_in), 
                      .pld_pma_tx_qpi_pulldn(pld_pma_tx_qpi_pulldn),
                      .pld_pma_tx_qpi_pullup(pld_pma_tx_qpi_pullup),
                      .pld_pma_rx_qpi_pullup(pld_pma_rx_qpi_pullup),
    
    // PLD DCM input
                      .pld_rx_clk1_dcm(pld_rx_clk1_dcm),
                      .pld_tx_clk1_dcm(pld_rx_clk1_dcm),
                      .pld_tx_clk2_dcm(pld_rx_clk2_dcm),
    
    // uC AVMM
    
    // DFT input
                      .dft_adpt_aibiobsr_fastclkn(1'b1),
                      .adapter_scan_rst_n(1'b1),
                      .adapter_scan_mode_n(1'b1),
                      .adapter_scan_shift_n(1'b1),
                      .adapter_scan_shift_clk(1'b0),
                      .adapter_scan_user_clk0(adapter_scan_user_clk0),         // 125MHz
                      .adapter_scan_user_clk1(adapter_scan_user_clk1),         // 250MHz
                      .adapter_scan_user_clk2(adapter_scan_user_clk2),         // 500MHz
                      .adapter_scan_user_clk3(adapter_scan_user_clk3),         // 1GHz
                      .adapter_clk_sel_n(1'b0),
                      .adapter_occ_enable(1'b0),
                      .adapter_global_pipe_se(1'b1),
                      .adapter_config_scan_in(4'h0),
                      .adapter_scan_in_occ1(2'h0),
                      .adapter_scan_in_occ2(5'h0),
                      .adapter_scan_in_occ3(1'b0),
                      .adapter_scan_in_occ4(1'b0),
                      .adapter_scan_in_occ5(2'h0),
                      .adapter_scan_in_occ6(11'h0),
                      .adapter_scan_in_occ7(1'b0),
                      .adapter_scan_in_occ8(1'b0),
                      .adapter_scan_in_occ9(1'b0),
                      .adapter_scan_in_occ10(1'b0),
                      .adapter_scan_in_occ11(1'b0),
                      .adapter_scan_in_occ12(1'b0),
                      .adapter_scan_in_occ13(1'b0),
                      .adapter_scan_in_occ14(1'b0),
                      .adapter_scan_in_occ15(1'b0),
                      .adapter_scan_in_occ16(1'b0),
                      .adapter_scan_in_occ17(1'b0),
                      .adapter_scan_in_occ18(2'h0),
                      .adapter_scan_in_occ19(1'h0),
                      .adapter_scan_in_occ20(1'h0),
                      .adapter_scan_in_occ21(2'h0),
                      .adapter_non_occ_scan_in(1'b0),
                      .adapter_occ_scan_in(1'b0),
                      .dft_fabric_iaibdftcore2dll(3'h0),
    
    
    // DFT output
                      .adapter_config_scan_out(),
                      .adapter_scan_out_occ1(),
                      .adapter_scan_out_occ2(),
                      .adapter_scan_out_occ3(),
                      .adapter_scan_out_occ4(),
                      .adapter_scan_out_occ5(),
                      .adapter_scan_out_occ6(),
                      .adapter_scan_out_occ7(),
                      .adapter_scan_out_occ8(),
                      .adapter_scan_out_occ9(),
                      .adapter_scan_out_occ10(),
                      .adapter_scan_out_occ11(),
                      .adapter_scan_out_occ12(),
                      .adapter_scan_out_occ13(),
                      .adapter_scan_out_occ14(),
                      .adapter_scan_out_occ15(),
                      .adapter_scan_out_occ16(),
                      .adapter_scan_out_occ17(),
                      .adapter_scan_out_occ18(),
                      .adapter_scan_out_occ19(),
                      .adapter_scan_out_occ20(),
                      .adapter_scan_out_occ21(),
                      .adapter_non_occ_scan_out(),
                      .adapter_occ_scan_out(),
                      .dft_fabric_oaibdftdll2core(),
    
    // Adapter output
                      .bond_rx_asn_ds_out_fifo_hold(),
                      .bond_rx_asn_us_out_fifo_hold(),
                      .bond_rx_fifo_ds_out_rden(),
                      .bond_rx_fifo_ds_out_wren(),
                      .bond_rx_fifo_us_out_rden(),
                      .bond_rx_fifo_us_out_wren(),
                      .bond_rx_hrdrst_ds_out_fabric_rx_dll_lock(),
                      .bond_rx_hrdrst_us_out_fabric_rx_dll_lock(),
                      .bond_rx_hrdrst_ds_out_fabric_rx_dll_lock_req(),
                      .bond_rx_hrdrst_us_out_fabric_rx_dll_lock_req(),
                      .bond_tx_fifo_ds_out_dv(),
                      .bond_tx_fifo_ds_out_rden(),
                      .bond_tx_fifo_ds_out_wren(),
                      .bond_tx_fifo_us_out_dv(),
                      .bond_tx_fifo_us_out_rden(),
                      .bond_tx_fifo_us_out_wren(),
                      .bond_tx_hrdrst_ds_out_fabric_tx_dcd_cal_done(),
                      .bond_tx_hrdrst_us_out_fabric_tx_dcd_cal_done(),
                      .bond_tx_hrdrst_ds_out_fabric_tx_dcd_cal_req(),
                      .bond_tx_hrdrst_us_out_fabric_tx_dcd_cal_req(),
    // Config output
                      .csr_clk_out(),
                      .csr_out(),
                      .csr_pipe_out(),
                      .csr_rdy_dly_out(),
                      .csr_rdy_out(),
                      .nfrzdrv_out(),
                      .usermode_out(),
    // PLD  output
                      .hip_aib_fsr_out(),
                      .hip_aib_ssr_out(),
                      .hip_avmm_readdata(),
                      .hip_avmm_readdatavalid(),
                      .hip_avmm_writedone(),
                      .hip_avmm_reserved_out(),
                      .pld_10g_krfec_rx_blk_lock(),
                      .pld_10g_krfec_rx_diag_data_status(),
                      .pld_10g_krfec_rx_frame(),
                      .pld_10g_krfec_tx_frame(),
                      .pld_krfec_tx_alignment(),
                      .pld_10g_rx_crc32_err(),
                      .pld_rx_fabric_fifo_insert(),
                      .pld_rx_fabric_fifo_del(),

                      .pld_10g_rx_frame_lock(),
                      .pld_10g_rx_hi_ber(),
                      .pld_10g_tx_burst_en_exe(),
                      .pld_8g_a1a2_k1k2_flag(),
                      .pld_8g_empty_rmf(),
                      .pld_8g_full_rmf(),
                      .pld_8g_rxelecidle(),
                      .pld_8g_signal_detect_out(),
                      .pld_8g_wa_boundary(),
                      .pld_avmm1_busy(),
                      .pld_avmm1_cmdfifo_wr_full(),
                      .pld_avmm1_cmdfifo_wr_pfull(),
                      .pld_avmm1_readdata(),
                      .pld_avmm1_readdatavalid(),
                      .pld_avmm1_reserved_out(),
                      .pld_avmm2_busy(),
                      .pld_avmm2_cmdfifo_wr_full(),
                      .pld_avmm2_cmdfifo_wr_pfull(),
                      .pld_avmm2_readdata(),
                      .pld_avmm2_readdatavalid(),
                      .pld_avmm2_reserved_out(),
                      .pld_chnl_cal_done(),
                      .pld_fpll_shared_direct_async_out(),
                      .pld_fpll_shared_direct_async_out_hioint(),
                      .pld_fpll_shared_direct_async_out_dcm(),
                      .pld_fsr_load(),
                      .pld_pcs_rx_clk_out1_hioint(),
                      .pld_pcs_rx_clk_out2_hioint(),
                      .pld_pcs_tx_clk_out1_hioint(),
                      .pld_pcs_tx_clk_out2_hioint(),
                      .pld_pll_cal_done(),
                      .pld_pma_adapt_done(),
                      .pld_pma_fpll_clk0bad(),
                      .pld_pma_fpll_clk1bad(),
                      .pld_pma_fpll_clksel(),
                      .pld_pma_fpll_phase_done(),
                      .pld_pma_hclk_hioint(),
                      .pld_pma_internal_clk1_hioint(),
                      .pld_pma_internal_clk2_hioint(),
                      .pld_pma_pcie_sw_done(),
                      .pld_pma_pfdmode_lock(),
                      .pld_pma_reserved_in(),
                      .pld_pma_rx_detect_valid(),
                      .pld_pma_rx_found(),
                      .pld_pma_rxpll_lock(),
                      .pld_pma_signal_ok(),
                      .pld_pma_testbus(),
                      .pld_pmaif_mask_tx_pll(),
                      .pld_rx_fabric_align_done(),
                      .pld_rx_fabric_data_out(pld_rx_fabric_data_out),
                      .pld_rx_fabric_fifo_empty(),
                      .pld_rx_fabric_fifo_full(),
                      .pld_rx_fabric_fifo_latency_pulse(),
                      .pld_rx_fabric_fifo_pempty(),
                      .pld_rx_fabric_fifo_pfull(),
                      .pld_rx_hssi_fifo_empty(),
                      .pld_rx_hssi_fifo_full(),
                      .pld_rx_hssi_fifo_latency_pulse(),
                      .pld_rx_prbs_done(),
                      .pld_rx_prbs_err(),
                      .pld_ssr_load(),
                      .pld_test_data(),
                      .pld_tx_fabric_fifo_empty(),
                      .pld_tx_fabric_fifo_full(),
                      .pld_tx_fabric_fifo_latency_pulse(),
                      .pld_tx_fabric_fifo_pempty(),
                      .pld_tx_fabric_fifo_pfull(),
                      .pld_tx_hssi_align_done(),
                      .pld_tx_hssi_fifo_empty(),
                      .pld_tx_hssi_fifo_full(),
                      .pld_tx_hssi_fifo_latency_pulse(),
                      .pld_hssi_osc_transfer_en(),
                      .pld_hssi_rx_transfer_en(),
                      .pld_fabric_tx_transfer_en(),
                      .pld_aib_fabric_rx_dll_lock(),
                      .pld_aib_fabric_tx_dcd_cal_done(),
                      .pld_aib_hssi_rx_dcd_cal_done(),
                      .pld_aib_hssi_tx_dcd_cal_done(),
                      .pld_aib_hssi_tx_dll_lock(),
                      .pld_hssi_asn_dll_lock_en(),
                      .pld_fabric_asn_dll_lock_en(),	
                      .pld_tx_ssr_reserved_out(),
                      .pld_rx_ssr_reserved_out(),
                          
                          // PLD DCM output
                      .pld_pcs_rx_clk_out1_dcm(),
                      .pld_pcs_rx_clk_out2_dcm(),
                      .pld_pcs_tx_clk_out1_dcm(),
                      .pld_pcs_tx_clk_out2_dcm(),

    //JTAG input
                      .iatpg_pipeline_global_en(1'b1),
                      .iatpg_scan_clk_in0(1'b1),
                      .iatpg_scan_clk_in1(1'b1),
                      .iatpg_scan_in0(1'b0),
                      .iatpg_scan_in1(1'b0),
                      .iatpg_scan_shift_n(1'b1),
                      .iatpg_scan_mode_n(1'b1),
                      .iatpg_scan_rst_n(1'b1),
                      .ijtag_clkdr_in_chain(1'b0),
                      .ijtag_last_bs_in_chain(1'b0),
                      .ijtag_tx_scan_in_chain(1'b0),
                      .ired_directin_data_in_chain1(ired_directin_data_in_chain1),
                      .ired_directin_data_in_chain2(ired_directin_data_in_chain2),
                      .ired_irxen_in_chain1(ired_irxen_in_chain1),
                      .ired_irxen_in_chain2(ired_irxen_in_chain2),
                      .ired_shift_en_in_chain1(ired_shift_en_in_chain1),
                      .ired_shift_en_in_chain2(ired_shift_en_in_chain2),
                      .jtag_clksel(1'b0),
                      .jtag_intest(1'b0),
                      .jtag_mode_in(1'b0),
                      .jtag_rstb(1'b1),
                      .jtag_rstb_en(1'b0),
                      .jtag_tx_scanen_in(1'b0),
                      .jtag_weakpdn(1'b0),
                      .jtag_weakpu(1'b0),

    //Jtag output 
                      .jtag_clksel_out(),
                      .jtag_intest_out(),
                      .jtag_mode_out(),
                      .jtag_rstb_en_out(),
                      .jtag_rstb_out(),
                      .jtag_tx_scanen_out(),
                      .jtag_weakpdn_out(),
                      .jtag_weakpu_out(),
                      .oatpg_scan_out0(),
                      .oatpg_scan_out1(),
                      .ojtag_clkdr_out_chain(),
                      .ojtag_last_bs_out_chain(),
                      .ojtag_rx_scan_out_chain(),
                      .ored_directin_data_out0_chain1(),
                      .ored_directin_data_out0_chain2(),
                      .ored_rxen_out_chain1(),
                      .ored_rxen_out_chain2(),
                      .ored_shift_en_out_chain1(),
                      .ored_shift_en_out_chain2()
);
    

