module emib_ch_m2s1 (
	inout [95:0] s_aib,
	inout [101:0] m_aib

	);

wire tie_low = 1'b0;

  aliasv xaliasv101 (
	.PLUS(m_aib[101]),
	.MINUS()
  );


  aliasv xaliasv100 (
	.PLUS(m_aib[100]),
	.MINUS()
  );

  aliasv xaliasv99 (
	.PLUS(m_aib[99]),
	.MINUS()
  );

  aliasv xaliasv98 (
	.PLUS(m_aib[98]),
	.MINUS()
  );


  aliasv xaliasv97 (
	.PLUS(m_aib[97]),
	.MINUS()
  );

  aliasv xaliasv96 (
	.PLUS(m_aib[96]),
	.MINUS()
  );

  aliasv xaliasv95 (
	.PLUS(m_aib[95]),
	.MINUS()
  );

  aliasv xaliasv94 (
	.PLUS(m_aib[94]),
	.MINUS()
  );

  aliasv xaliasv93 (
	.PLUS(m_aib[93]),
	.MINUS()
  );

  aliasv xaliasv92 (
	.PLUS(m_aib[92]),
	.MINUS()
  );

  aliasv xaliasv91 (
	.PLUS(m_aib[91]),
	.MINUS()
  );

  aliasv xaliasv90 (
	.PLUS(m_aib[90]),
	.MINUS()
  );

  aliasv xaliasv89 (
	.PLUS(m_aib[89]),
	.MINUS()
  );

  aliasv xaliasv88 (
	.PLUS(m_aib[88]),
	.MINUS()
  );

  aliasv xaliasv87 (
	.PLUS(m_aib[87]),
	.MINUS()
  );

  aliasv xaliasv86 (
	.PLUS(m_aib[86]),
	.MINUS()
  );

  aliasv xaliasv85 (
	.PLUS(m_aib[85]),
	.MINUS()
  );

  aliasv xaliasv84 (
	.PLUS(m_aib[84]),
	.MINUS()
  );

  aliasv xaliasv83 (
	.PLUS(m_aib[83]),
	.MINUS()
  );

  aliasv xaliasv82 (
	.PLUS(m_aib[82]),
	.MINUS()
  );

  aliasv xaliasv81 (
	.PLUS(m_aib[81]),
	.MINUS(s_aib[38])
  );

  aliasv xaliasv80 (
	.PLUS(m_aib[80]),
	.MINUS(s_aib[39])
  );

  aliasv xaliasv79 (
	.PLUS(m_aib[79]),
	.MINUS(s_aib[36])
  );

  aliasv xaliasv78 (
	.PLUS(m_aib[78]),
	.MINUS(s_aib[37])
  );

  aliasv xaliasv77 (
	.PLUS(m_aib[77]),
	.MINUS(s_aib[34])
  );

  aliasv xaliasv76 (
	.PLUS(m_aib[76]),
	.MINUS(s_aib[35])
  );

  aliasv xaliasv75 (
	.PLUS(m_aib[75]),
	.MINUS(s_aib[32])
  );

  aliasv xaliasv74 (
	.PLUS(m_aib[74]),
	.MINUS(s_aib[33])
  );

  aliasv xaliasv73 (
	.PLUS(m_aib[73]),
	.MINUS(s_aib[30])
  );

  aliasv xaliasv72 (
	.PLUS(m_aib[72]),
	.MINUS(s_aib[31])
  );

  aliasv xaliasv71 (
	.PLUS(m_aib[71]),
	.MINUS(s_aib[43])
  );

  aliasv xaliasv70 (
	.PLUS(m_aib[70]),
	.MINUS(s_aib[42])
  );

  aliasv xaliasv69 (
	.PLUS(m_aib[69]),
	.MINUS(s_aib[28])
  );

  aliasv xaliasv68 (
	.PLUS(m_aib[68]),
	.MINUS(s_aib[29])
  );

  aliasv xaliasv67 (
	.PLUS(m_aib[67]),
	.MINUS(s_aib[26])
  );

  aliasv xaliasv66 (
	.PLUS(m_aib[66]),
	.MINUS(s_aib[27])
  );

  aliasv xaliasv65 (
	.PLUS(m_aib[65]),
	.MINUS(s_aib[24])
  );

  aliasv xaliasv64 (
	.PLUS(m_aib[64]),
	.MINUS(s_aib[25])
  );

  aliasv xaliasv63 (
	.PLUS(m_aib[63]),
	.MINUS(s_aib[22])
  );

  aliasv xaliasv62 (
	.PLUS(m_aib[62]),
	.MINUS(s_aib[23])
  );

  aliasv xaliasv61 (
	.PLUS(m_aib[61]),
	.MINUS(s_aib[20])
  );

  aliasv xaliasv60 (
	.PLUS(m_aib[60]),
	.MINUS(s_aib[21])
  );

  aliasv xaliasv59 (
	.PLUS(m_aib[59]),
	.MINUS(s_aib[57])
  );

  aliasv xaliasv58 (
	.PLUS(m_aib[58]),
	.MINUS(s_aib[59])
  );

  aliasv xaliasv57 (
	.PLUS(m_aib[57]),
	.MINUS(s_aib[83])
  );

  aliasv xaliasv56 (
	.PLUS(m_aib[56]),
	.MINUS(s_aib[82])
  );

  aliasv xaliasv55 (
	.PLUS(m_aib[55]),
	.MINUS(s_aib[93])
  );

  aliasv xaliasv54 (
	.PLUS(m_aib[54]),
	.MINUS(s_aib[92])
  );

  aliasv xaliasv53 (
	.PLUS(m_aib[53]),
	.MINUS(s_aib[44])
  );

  aliasv xaliasv52 (
	.PLUS(m_aib[52]),
	.MINUS(s_aib[65])
  );

  aliasv xaliasv51 (
	.PLUS(m_aib[51]),
	.MINUS()
  );

  aliasv xaliasv50 (
	.PLUS(m_aib[50]),
	.MINUS()
  );

  aliasv xaliasv49 (
	.PLUS(m_aib[49]),
	.MINUS(s_aib[56])
  );

  aliasv xaliasv48 (
	.PLUS(m_aib[48]),
	.MINUS(s_aib[49])
  );

  aliasv xaliasv47 (
	.PLUS(m_aib[47]),
	.MINUS(s_aib[94])
  );

  aliasv xaliasv46 (
	.PLUS(m_aib[46]),
	.MINUS(s_aib[95])
  );

  aliasv xaliasv45 (
	.PLUS(m_aib[45]),
	.MINUS(s_aib[84])
  );

  aliasv xaliasv44 (
	.PLUS(m_aib[44]),
	.MINUS(s_aib[85])
  );

  aliasv xaliasv43 (
	.PLUS(m_aib[43]),
	.MINUS(s_aib[86])
  );

  aliasv xaliasv42 (
	.PLUS(m_aib[42]),
	.MINUS(s_aib[87])
  );

  aliasv xaliasv41 (
	.PLUS(m_aib[41]),
	.MINUS(s_aib[1])
  );

  aliasv xaliasv40 (
	.PLUS(m_aib[40]),
	.MINUS(s_aib[0])
  );

  aliasv xaliasv39 (
	.PLUS(m_aib[39]),
	.MINUS(s_aib[3])
  );

  aliasv xaliasv38 (
	.PLUS(m_aib[38]),
	.MINUS(s_aib[2])
  );

  aliasv xaliasv37 (
	.PLUS(m_aib[37]),
	.MINUS(s_aib[5])
  );

  aliasv xaliasv36 (
	.PLUS(m_aib[36]),
	.MINUS(s_aib[4])
  );

  aliasv xaliasv35 (
	.PLUS(m_aib[35]),
	.MINUS(s_aib[7])
  );

  aliasv xaliasv34 (
	.PLUS(m_aib[34]),
	.MINUS(s_aib[6])
  );

  aliasv xaliasv33 (
	.PLUS(m_aib[33]),
	.MINUS(s_aib[9])
  );

  aliasv xaliasv32 (
	.PLUS(m_aib[32]),
	.MINUS(s_aib[8])
  );

  aliasv xaliasv31 (
	.PLUS(m_aib[31]),
	.MINUS(s_aib[40])
  );

  aliasv xaliasv30 (
	.PLUS(m_aib[30]),
	.MINUS(s_aib[41])
  );

  aliasv xaliasv29 (
	.PLUS(m_aib[29]),
	.MINUS(s_aib[11])
  );

  aliasv xaliasv28 (
	.PLUS(m_aib[28]),
	.MINUS(s_aib[10])
  );

  aliasv xaliasv27 (
	.PLUS(m_aib[27]),
	.MINUS(s_aib[13])
  );

  aliasv xaliasv26 (
	.PLUS(m_aib[26]),
	.MINUS(s_aib[12])
  );

  aliasv xaliasv25 (
	.PLUS(m_aib[25]),
	.MINUS(s_aib[15])
  );

  aliasv xaliasv24 (
	.PLUS(m_aib[24]),
	.MINUS(s_aib[14])
  );

  aliasv xaliasv23 (
	.PLUS(m_aib[23]),
	.MINUS(s_aib[17])
  );

  aliasv xaliasv22 (
	.PLUS(m_aib[22]),
	.MINUS(s_aib[16])
  );

  aliasv xaliasv21 (
	.PLUS(m_aib[21]),
	.MINUS(s_aib[19])
  );

  aliasv xaliasv20 (
	.PLUS(m_aib[20]),
	.MINUS(s_aib[18])
  );

  aliasv xaliasv19 (
	.PLUS(m_aib[19]),
	.MINUS()
  );

  aliasv xaliasv18 (
	.PLUS(m_aib[18]),
	.MINUS()
  );

  aliasv xaliasv17 (
	.PLUS(m_aib[17]),
	.MINUS()
  );

  aliasv xaliasv16 (
	.PLUS(m_aib[16]),
	.MINUS()
  );

  aliasv xaliasv15 (
	.PLUS(m_aib[15]),
	.MINUS()
  );

  aliasv xaliasv14 (
	.PLUS(m_aib[14]),
	.MINUS()
  );

  aliasv xaliasv13 (
	.PLUS(m_aib[13]),
	.MINUS()
  );

  aliasv xaliasv12 (
	.PLUS(m_aib[12]),
	.MINUS()
  );

  aliasv xaliasv11 (
	.PLUS(m_aib[11]),
	.MINUS()
  );

  aliasv xaliasv10 (
	.PLUS(m_aib[10]),
	.MINUS()
  );

  aliasv xaliasv9 (
	.PLUS(m_aib[9]),
	.MINUS()
  );

  aliasv xaliasv8 (
	.PLUS(m_aib[8]),
	.MINUS()
  );

  aliasv xaliasv7 (
	.PLUS(m_aib[7]),
	.MINUS()
  );

  aliasv xaliasv6 (
	.PLUS(m_aib[6]),
	.MINUS()
  );

  aliasv xaliasv5 (
	.PLUS(m_aib[5]),
	.MINUS()
  );

  aliasv xaliasv4 (
	.PLUS(m_aib[4]),
	.MINUS()
  );

  aliasv xaliasv3 (
	.PLUS(m_aib[3]),
	.MINUS()
  );

  aliasv xaliasv2 (
	.PLUS(m_aib[2]),
	.MINUS()
  );

  aliasv xaliasv1 (
	.PLUS(m_aib[1]),
	.MINUS()
  );

  aliasv xaliasv0 (
	.PLUS(m_aib[0]),
	.MINUS()
  );

//Unused pin of Slave MAIB
  aliasv xalias_sl45 (
        .PLUS(),
        .MINUS(s_aib[45])
  );

  aliasv xalias_sl58 (
        .PLUS(),
        .MINUS(s_aib[58])
  );


  aliasv xalias_sl61 (
        .PLUS(),
        .MINUS(s_aib[61])
  );

  aliasv xalias_sl63 (
        .PLUS(),
        .MINUS(s_aib[63])
  );

  aliasv xalias_sl64 (
        .PLUS(),
        .MINUS(s_aib[64])
  );

  aliasv xalias_sl67 (
        .PLUS(),
        .MINUS(s_aib[67])
  );

  aliasv xalias_sl73 (
        .PLUS(),
        .MINUS(s_aib[73])
  );

  aliasv xalias_sl74 (
        .PLUS(),
        .MINUS(s_aib[74])
  );

  aliasv xalias_sl78 (
        .PLUS(),
        .MINUS(s_aib[78])
  );

  aliasv xalias_sl79 (
        .PLUS(),
        .MINUS(s_aib[79])
  );

  aliasv xalias_sl80 (
        .PLUS(),
        .MINUS(s_aib[80])
  );

  aliasv xalias_sl81 (
        .PLUS(),
        .MINUS(s_aib[81])
  );

  aliasv xalias_sl88 (
        .PLUS(),
        .MINUS(s_aib[88])
  );

  aliasv xalias_sl89 (
        .PLUS(),
        .MINUS(s_aib[89])
  );

  aliasv xalias_sl47 (
        .PLUS(tie_low),
        .MINUS(s_aib[47])
  );

  aliasv xalias_sl46 (
        .PLUS(tie_low),
        .MINUS(s_aib[46])
  );

  aliasv xalias_sl48 (
        .PLUS(tie_low),
        .MINUS(s_aib[48])
  );


  aliasv xalias_sl50 (
        .PLUS(tie_low),
        .MINUS(s_aib[50])
  );

  aliasv xalias_sl51 (
        .PLUS(tie_low),
        .MINUS(s_aib[51])
  );

  aliasv xalias_sl52 (
        .PLUS(tie_low),
        .MINUS(s_aib[52])
  );

  aliasv xalias_sl53 (
        .PLUS(tie_low),
        .MINUS(s_aib[53])
  );

  aliasv xalias_sl54 (
        .PLUS(tie_low),
        .MINUS(s_aib[54])
  );

  aliasv xalias_sl55 (
        .PLUS(tie_low),
        .MINUS(s_aib[55])
  );

  aliasv xalias_sl60 (
        .PLUS(tie_low),
        .MINUS(s_aib[60])
  );

  aliasv xalias_sl62 (
        .PLUS(tie_low),
        .MINUS(s_aib[62])
  );


  aliasv xalias_sl66 (
        .PLUS(tie_low),
        .MINUS(s_aib[66])
  );


  aliasv xalias_sl68 (
        .PLUS(tie_low),
        .MINUS(s_aib[68])
  );


  aliasv xalias_sl69 (
        .PLUS(tie_low),
        .MINUS(s_aib[69])
  );

  aliasv xalias_sl70 (
        .PLUS(tie_low),
        .MINUS(s_aib[70])
  );

  aliasv xalias_sl71 (
        .PLUS(tie_low),
        .MINUS(s_aib[71])
  );

  aliasv xalias_sl72 (
        .PLUS(),
        .MINUS(s_aib[72])
  );

  aliasv xalias_sl75 (
        .PLUS(tie_low),
        .MINUS(s_aib[75])
  );

  aliasv xalias_sl76 (
        .PLUS(tie_low),
        .MINUS(s_aib[76])
  );

  aliasv xalias_sl77 (
        .PLUS(tie_low),
        .MINUS(s_aib[77])
  );

  aliasv xalias_sl90 (
        .PLUS(tie_low),
        .MINUS(s_aib[90])
  );

  aliasv xalias_sl91 (
        .PLUS(tie_low),
        .MINUS(s_aib[91])
  );
endmodule
