// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. All rights reserved
module aibnd_aliasd ( PLUS, MINUS );

	input   PLUS;
	output  MINUS;

	assign MINUS = PLUS;

endmodule





