// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. 
// *****************************************************************************
// *****************************************************************************
//  Copyright © 2016 Altera Corporation.  
// *****************************************************************************
//  Module Name :  c3lib_ecc_enc_d80_c88
//  Date        :  Mon May 16 22:06:38 2016
//  Description :  ECC encoder (based on the standard Extended Hamming Code
//                 scheme). Code generated by ecc_gen.pl script (command line
//                 options used: -num_data_bits 80).
// *****************************************************************************

module c3lib_ecc_enc_d80_c88(

  input  logic[ 79 : 0 ]	i_data,
  output logic[ 87 : 0 ]	o_code

);

assign o_code[ 0 ] = o_code[ 1 ] ^ o_code[ 2 ] ^ o_code[ 3 ] ^ o_code[ 4 ] ^ o_code[ 5 ] ^ o_code[ 6 ] ^ o_code[ 7 ] ^ o_code[ 8 ] ^ o_code[ 9 ] ^ o_code[ 10 ] ^ o_code[ 11 ] ^ o_code[ 12 ] ^ o_code[ 13 ] ^ o_code[ 14 ] ^ o_code[ 15 ] ^ o_code[ 16 ] ^ o_code[ 17 ] ^ o_code[ 18 ] ^ o_code[ 19 ] ^ o_code[ 20 ] ^ o_code[ 21 ] ^ o_code[ 22 ] ^ o_code[ 23 ] ^ o_code[ 24 ] ^ o_code[ 25 ] ^ o_code[ 26 ] ^ o_code[ 27 ] ^ o_code[ 28 ] ^ o_code[ 29 ] ^ o_code[ 30 ] ^ o_code[ 31 ] ^ o_code[ 32 ] ^ o_code[ 33 ] ^ o_code[ 34 ] ^ o_code[ 35 ] ^ o_code[ 36 ] ^ o_code[ 37 ] ^ o_code[ 38 ] ^ o_code[ 39 ] ^ o_code[ 40 ] ^ o_code[ 41 ] ^ o_code[ 42 ] ^ o_code[ 43 ] ^ o_code[ 44 ] ^ o_code[ 45 ] ^ o_code[ 46 ] ^ o_code[ 47 ] ^ o_code[ 48 ] ^ o_code[ 49 ] ^ o_code[ 50 ] ^ o_code[ 51 ] ^ o_code[ 52 ] ^ o_code[ 53 ] ^ o_code[ 54 ] ^ o_code[ 55 ] ^ o_code[ 56 ] ^ o_code[ 57 ] ^ o_code[ 58 ] ^ o_code[ 59 ] ^ o_code[ 60 ] ^ o_code[ 61 ] ^ o_code[ 62 ] ^ o_code[ 63 ] ^ o_code[ 64 ] ^ o_code[ 65 ] ^ o_code[ 66 ] ^ o_code[ 67 ] ^ o_code[ 68 ] ^ o_code[ 69 ] ^ o_code[ 70 ] ^ o_code[ 71 ] ^ o_code[ 72 ] ^ o_code[ 73 ] ^ o_code[ 74 ] ^ o_code[ 75 ] ^ o_code[ 76 ] ^ o_code[ 77 ] ^ o_code[ 78 ] ^ o_code[ 79 ] ^ o_code[ 80 ] ^ o_code[ 81 ] ^ o_code[ 82 ] ^ o_code[ 83 ] ^ o_code[ 84 ] ^ o_code[ 85 ] ^ o_code[ 86 ] ^ o_code[ 87 ];
assign o_code[ 1 ] = o_code[ 3 ] ^ o_code[ 5 ] ^ o_code[ 7 ] ^ o_code[ 9 ] ^ o_code[ 11 ] ^ o_code[ 13 ] ^ o_code[ 15 ] ^ o_code[ 17 ] ^ o_code[ 19 ] ^ o_code[ 21 ] ^ o_code[ 23 ] ^ o_code[ 25 ] ^ o_code[ 27 ] ^ o_code[ 29 ] ^ o_code[ 31 ] ^ o_code[ 33 ] ^ o_code[ 35 ] ^ o_code[ 37 ] ^ o_code[ 39 ] ^ o_code[ 41 ] ^ o_code[ 43 ] ^ o_code[ 45 ] ^ o_code[ 47 ] ^ o_code[ 49 ] ^ o_code[ 51 ] ^ o_code[ 53 ] ^ o_code[ 55 ] ^ o_code[ 57 ] ^ o_code[ 59 ] ^ o_code[ 61 ] ^ o_code[ 63 ] ^ o_code[ 65 ] ^ o_code[ 67 ] ^ o_code[ 69 ] ^ o_code[ 71 ] ^ o_code[ 73 ] ^ o_code[ 75 ] ^ o_code[ 77 ] ^ o_code[ 79 ] ^ o_code[ 81 ] ^ o_code[ 83 ] ^ o_code[ 85 ] ^ o_code[ 87 ];
assign o_code[ 2 ] = o_code[ 3 ] ^ o_code[ 6 ] ^ o_code[ 7 ] ^ o_code[ 10 ] ^ o_code[ 11 ] ^ o_code[ 14 ] ^ o_code[ 15 ] ^ o_code[ 18 ] ^ o_code[ 19 ] ^ o_code[ 22 ] ^ o_code[ 23 ] ^ o_code[ 26 ] ^ o_code[ 27 ] ^ o_code[ 30 ] ^ o_code[ 31 ] ^ o_code[ 34 ] ^ o_code[ 35 ] ^ o_code[ 38 ] ^ o_code[ 39 ] ^ o_code[ 42 ] ^ o_code[ 43 ] ^ o_code[ 46 ] ^ o_code[ 47 ] ^ o_code[ 50 ] ^ o_code[ 51 ] ^ o_code[ 54 ] ^ o_code[ 55 ] ^ o_code[ 58 ] ^ o_code[ 59 ] ^ o_code[ 62 ] ^ o_code[ 63 ] ^ o_code[ 66 ] ^ o_code[ 67 ] ^ o_code[ 70 ] ^ o_code[ 71 ] ^ o_code[ 74 ] ^ o_code[ 75 ] ^ o_code[ 78 ] ^ o_code[ 79 ] ^ o_code[ 82 ] ^ o_code[ 83 ] ^ o_code[ 86 ] ^ o_code[ 87 ];
assign o_code[ 3 ] = i_data[ 0 ];
assign o_code[ 4 ] = o_code[ 5 ] ^ o_code[ 6 ] ^ o_code[ 7 ] ^ o_code[ 12 ] ^ o_code[ 13 ] ^ o_code[ 14 ] ^ o_code[ 15 ] ^ o_code[ 20 ] ^ o_code[ 21 ] ^ o_code[ 22 ] ^ o_code[ 23 ] ^ o_code[ 28 ] ^ o_code[ 29 ] ^ o_code[ 30 ] ^ o_code[ 31 ] ^ o_code[ 36 ] ^ o_code[ 37 ] ^ o_code[ 38 ] ^ o_code[ 39 ] ^ o_code[ 44 ] ^ o_code[ 45 ] ^ o_code[ 46 ] ^ o_code[ 47 ] ^ o_code[ 52 ] ^ o_code[ 53 ] ^ o_code[ 54 ] ^ o_code[ 55 ] ^ o_code[ 60 ] ^ o_code[ 61 ] ^ o_code[ 62 ] ^ o_code[ 63 ] ^ o_code[ 68 ] ^ o_code[ 69 ] ^ o_code[ 70 ] ^ o_code[ 71 ] ^ o_code[ 76 ] ^ o_code[ 77 ] ^ o_code[ 78 ] ^ o_code[ 79 ] ^ o_code[ 84 ] ^ o_code[ 85 ] ^ o_code[ 86 ] ^ o_code[ 87 ];
assign o_code[ 5 ] = i_data[ 1 ];
assign o_code[ 6 ] = i_data[ 2 ];
assign o_code[ 7 ] = i_data[ 3 ];
assign o_code[ 8 ] = o_code[ 9 ] ^ o_code[ 10 ] ^ o_code[ 11 ] ^ o_code[ 12 ] ^ o_code[ 13 ] ^ o_code[ 14 ] ^ o_code[ 15 ] ^ o_code[ 24 ] ^ o_code[ 25 ] ^ o_code[ 26 ] ^ o_code[ 27 ] ^ o_code[ 28 ] ^ o_code[ 29 ] ^ o_code[ 30 ] ^ o_code[ 31 ] ^ o_code[ 40 ] ^ o_code[ 41 ] ^ o_code[ 42 ] ^ o_code[ 43 ] ^ o_code[ 44 ] ^ o_code[ 45 ] ^ o_code[ 46 ] ^ o_code[ 47 ] ^ o_code[ 56 ] ^ o_code[ 57 ] ^ o_code[ 58 ] ^ o_code[ 59 ] ^ o_code[ 60 ] ^ o_code[ 61 ] ^ o_code[ 62 ] ^ o_code[ 63 ] ^ o_code[ 72 ] ^ o_code[ 73 ] ^ o_code[ 74 ] ^ o_code[ 75 ] ^ o_code[ 76 ] ^ o_code[ 77 ] ^ o_code[ 78 ] ^ o_code[ 79 ];
assign o_code[ 9 ] = i_data[ 4 ];
assign o_code[ 10 ] = i_data[ 5 ];
assign o_code[ 11 ] = i_data[ 6 ];
assign o_code[ 12 ] = i_data[ 7 ];
assign o_code[ 13 ] = i_data[ 8 ];
assign o_code[ 14 ] = i_data[ 9 ];
assign o_code[ 15 ] = i_data[ 10 ];
assign o_code[ 16 ] = o_code[ 17 ] ^ o_code[ 18 ] ^ o_code[ 19 ] ^ o_code[ 20 ] ^ o_code[ 21 ] ^ o_code[ 22 ] ^ o_code[ 23 ] ^ o_code[ 24 ] ^ o_code[ 25 ] ^ o_code[ 26 ] ^ o_code[ 27 ] ^ o_code[ 28 ] ^ o_code[ 29 ] ^ o_code[ 30 ] ^ o_code[ 31 ] ^ o_code[ 48 ] ^ o_code[ 49 ] ^ o_code[ 50 ] ^ o_code[ 51 ] ^ o_code[ 52 ] ^ o_code[ 53 ] ^ o_code[ 54 ] ^ o_code[ 55 ] ^ o_code[ 56 ] ^ o_code[ 57 ] ^ o_code[ 58 ] ^ o_code[ 59 ] ^ o_code[ 60 ] ^ o_code[ 61 ] ^ o_code[ 62 ] ^ o_code[ 63 ] ^ o_code[ 80 ] ^ o_code[ 81 ] ^ o_code[ 82 ] ^ o_code[ 83 ] ^ o_code[ 84 ] ^ o_code[ 85 ] ^ o_code[ 86 ] ^ o_code[ 87 ];
assign o_code[ 17 ] = i_data[ 11 ];
assign o_code[ 18 ] = i_data[ 12 ];
assign o_code[ 19 ] = i_data[ 13 ];
assign o_code[ 20 ] = i_data[ 14 ];
assign o_code[ 21 ] = i_data[ 15 ];
assign o_code[ 22 ] = i_data[ 16 ];
assign o_code[ 23 ] = i_data[ 17 ];
assign o_code[ 24 ] = i_data[ 18 ];
assign o_code[ 25 ] = i_data[ 19 ];
assign o_code[ 26 ] = i_data[ 20 ];
assign o_code[ 27 ] = i_data[ 21 ];
assign o_code[ 28 ] = i_data[ 22 ];
assign o_code[ 29 ] = i_data[ 23 ];
assign o_code[ 30 ] = i_data[ 24 ];
assign o_code[ 31 ] = i_data[ 25 ];
assign o_code[ 32 ] = o_code[ 33 ] ^ o_code[ 34 ] ^ o_code[ 35 ] ^ o_code[ 36 ] ^ o_code[ 37 ] ^ o_code[ 38 ] ^ o_code[ 39 ] ^ o_code[ 40 ] ^ o_code[ 41 ] ^ o_code[ 42 ] ^ o_code[ 43 ] ^ o_code[ 44 ] ^ o_code[ 45 ] ^ o_code[ 46 ] ^ o_code[ 47 ] ^ o_code[ 48 ] ^ o_code[ 49 ] ^ o_code[ 50 ] ^ o_code[ 51 ] ^ o_code[ 52 ] ^ o_code[ 53 ] ^ o_code[ 54 ] ^ o_code[ 55 ] ^ o_code[ 56 ] ^ o_code[ 57 ] ^ o_code[ 58 ] ^ o_code[ 59 ] ^ o_code[ 60 ] ^ o_code[ 61 ] ^ o_code[ 62 ] ^ o_code[ 63 ];
assign o_code[ 33 ] = i_data[ 26 ];
assign o_code[ 34 ] = i_data[ 27 ];
assign o_code[ 35 ] = i_data[ 28 ];
assign o_code[ 36 ] = i_data[ 29 ];
assign o_code[ 37 ] = i_data[ 30 ];
assign o_code[ 38 ] = i_data[ 31 ];
assign o_code[ 39 ] = i_data[ 32 ];
assign o_code[ 40 ] = i_data[ 33 ];
assign o_code[ 41 ] = i_data[ 34 ];
assign o_code[ 42 ] = i_data[ 35 ];
assign o_code[ 43 ] = i_data[ 36 ];
assign o_code[ 44 ] = i_data[ 37 ];
assign o_code[ 45 ] = i_data[ 38 ];
assign o_code[ 46 ] = i_data[ 39 ];
assign o_code[ 47 ] = i_data[ 40 ];
assign o_code[ 48 ] = i_data[ 41 ];
assign o_code[ 49 ] = i_data[ 42 ];
assign o_code[ 50 ] = i_data[ 43 ];
assign o_code[ 51 ] = i_data[ 44 ];
assign o_code[ 52 ] = i_data[ 45 ];
assign o_code[ 53 ] = i_data[ 46 ];
assign o_code[ 54 ] = i_data[ 47 ];
assign o_code[ 55 ] = i_data[ 48 ];
assign o_code[ 56 ] = i_data[ 49 ];
assign o_code[ 57 ] = i_data[ 50 ];
assign o_code[ 58 ] = i_data[ 51 ];
assign o_code[ 59 ] = i_data[ 52 ];
assign o_code[ 60 ] = i_data[ 53 ];
assign o_code[ 61 ] = i_data[ 54 ];
assign o_code[ 62 ] = i_data[ 55 ];
assign o_code[ 63 ] = i_data[ 56 ];
assign o_code[ 64 ] = o_code[ 65 ] ^ o_code[ 66 ] ^ o_code[ 67 ] ^ o_code[ 68 ] ^ o_code[ 69 ] ^ o_code[ 70 ] ^ o_code[ 71 ] ^ o_code[ 72 ] ^ o_code[ 73 ] ^ o_code[ 74 ] ^ o_code[ 75 ] ^ o_code[ 76 ] ^ o_code[ 77 ] ^ o_code[ 78 ] ^ o_code[ 79 ] ^ o_code[ 80 ] ^ o_code[ 81 ] ^ o_code[ 82 ] ^ o_code[ 83 ] ^ o_code[ 84 ] ^ o_code[ 85 ] ^ o_code[ 86 ] ^ o_code[ 87 ];
assign o_code[ 65 ] = i_data[ 57 ];
assign o_code[ 66 ] = i_data[ 58 ];
assign o_code[ 67 ] = i_data[ 59 ];
assign o_code[ 68 ] = i_data[ 60 ];
assign o_code[ 69 ] = i_data[ 61 ];
assign o_code[ 70 ] = i_data[ 62 ];
assign o_code[ 71 ] = i_data[ 63 ];
assign o_code[ 72 ] = i_data[ 64 ];
assign o_code[ 73 ] = i_data[ 65 ];
assign o_code[ 74 ] = i_data[ 66 ];
assign o_code[ 75 ] = i_data[ 67 ];
assign o_code[ 76 ] = i_data[ 68 ];
assign o_code[ 77 ] = i_data[ 69 ];
assign o_code[ 78 ] = i_data[ 70 ];
assign o_code[ 79 ] = i_data[ 71 ];
assign o_code[ 80 ] = i_data[ 72 ];
assign o_code[ 81 ] = i_data[ 73 ];
assign o_code[ 82 ] = i_data[ 74 ];
assign o_code[ 83 ] = i_data[ 75 ];
assign o_code[ 84 ] = i_data[ 76 ];
assign o_code[ 85 ] = i_data[ 77 ];
assign o_code[ 86 ] = i_data[ 78 ];
assign o_code[ 87 ] = i_data[ 79 ];

endmodule

