module emib_ch (
	inout s_aib95,
	inout aib95,
	inout s_aib94,
	inout aib94,
	inout s_aib93,
	inout aib93,
	inout s_aib92,
	inout aib92,
	inout s_aib91,
	inout aib91,
	inout s_aib90,
	inout aib90,
	inout s_aib89,
	inout aib89,
	inout s_aib88,
	inout aib88,
	inout s_aib87,
	inout aib87,
	inout s_aib86,
	inout aib86,
	inout s_aib85,
	inout aib85,
	inout s_aib84,
	inout aib84,
	inout s_aib83,
	inout aib83,
	inout s_aib82,
	inout aib82,
	inout s_aib81,
	inout aib81,
	inout s_aib80,
	inout aib80,
	inout s_aib79,
	inout aib79,
	inout s_aib78,
	inout aib78,
	inout s_aib77,
	inout aib77,
	inout s_aib76,
	inout aib76,
	inout s_aib75,
	inout aib75,
	inout s_aib74,
	inout aib74,
	inout s_aib73,
	inout aib73,
	inout s_aib72,
	inout aib72,
	inout s_aib71,
	inout aib71,
	inout s_aib70,
	inout aib70,
	inout s_aib69,
	inout aib69,
	inout s_aib68,
	inout aib68,
	inout s_aib67,
	inout aib67,
	inout s_aib66,
	inout aib66,
	inout s_aib65,
	inout aib65,
	inout s_aib64,
	inout aib64,
	inout s_aib63,
	inout aib63,
	inout s_aib62,
	inout aib62,
	inout s_aib61,
	inout aib61,
	inout s_aib60,
	inout aib60,
	inout s_aib59,
	inout aib59,
	inout s_aib58,
	inout aib58,
	inout s_aib57,
	inout aib57,
	inout s_aib56,
	inout aib56,
	inout s_aib55,
	inout aib55,
	inout s_aib54,
	inout aib54,
	inout s_aib53,
	inout aib53,
	inout s_aib52,
	inout aib52,
	inout s_aib51,
	inout aib51,
	inout s_aib50,
	inout aib50,
	inout s_aib49,
	inout aib49,
	inout s_aib48,
	inout aib48,
	inout s_aib47,
	inout aib47,
	inout s_aib46,
	inout aib46,
	inout s_aib45,
	inout aib45,
	inout s_aib44,
	inout aib44,
	inout s_aib43,
	inout aib43,
	inout s_aib42,
	inout aib42,
	inout s_aib41,
	inout aib41,
	inout s_aib40,
	inout aib40,
	inout s_aib39,
	inout aib39,
	inout s_aib38,
	inout aib38,
	inout s_aib37,
	inout aib37,
	inout s_aib36,
	inout aib36,
	inout s_aib35,
	inout aib35,
	inout s_aib34,
	inout aib34,
	inout s_aib33,
	inout aib33,
	inout s_aib32,
	inout aib32,
	inout s_aib31,
	inout aib31,
	inout s_aib30,
	inout aib30,
	inout s_aib29,
	inout aib29,
	inout s_aib28,
	inout aib28,
	inout s_aib27,
	inout aib27,
	inout s_aib26,
	inout aib26,
	inout s_aib25,
	inout aib25,
	inout s_aib24,
	inout aib24,
	inout s_aib23,
	inout aib23,
	inout s_aib22,
	inout aib22,
	inout s_aib21,
	inout aib21,
	inout s_aib20,
	inout aib20,
	inout s_aib19,
	inout aib19,
	inout s_aib18,
	inout aib18,
	inout s_aib17,
	inout aib17,
	inout s_aib16,
	inout aib16,
	inout s_aib15,
	inout aib15,
	inout s_aib14,
	inout aib14,
	inout s_aib13,
	inout aib13,
	inout s_aib12,
	inout aib12,
	inout s_aib11,
	inout aib11,
	inout s_aib10,
	inout aib10,
	inout s_aib9,
	inout aib9,
	inout s_aib8,
	inout aib8,
	inout s_aib7,
	inout aib7,
	inout s_aib6,
	inout aib6,
	inout s_aib5,
	inout aib5,
	inout s_aib4,
	inout aib4,
	inout s_aib3,
	inout aib3,
	inout s_aib2,
	inout aib2,
	inout s_aib1,
	inout aib1,
	inout s_aib0,
	inout aib0

	);
  aliasv xaliasv95 (
	.PLUS(s_aib95),
	.MINUS(aib95)
  );

  aliasv xaliasv94 (
	.PLUS(s_aib94),
	.MINUS(aib94)
  );

  aliasv xaliasv93 (
	.PLUS(s_aib93),
	.MINUS(aib93)
  );

  aliasv xaliasv92 (
	.PLUS(s_aib92),
	.MINUS(aib92)
  );

  aliasv xaliasv91 (
	.PLUS(s_aib91),
	.MINUS(aib91)
  );

  aliasv xaliasv90 (
	.PLUS(s_aib90),
	.MINUS(aib90)
  );

  aliasv xaliasv89 (
	.PLUS(s_aib89),
	.MINUS(aib89)
  );

  aliasv xaliasv88 (
	.PLUS(s_aib88),
	.MINUS(aib88)
  );

  aliasv xaliasv87 (
	.PLUS(s_aib87),
	.MINUS(aib87)
  );

  aliasv xaliasv86 (
	.PLUS(s_aib86),
	.MINUS(aib86)
  );

  aliasv xaliasv85 (
	.PLUS(s_aib85),
	.MINUS(aib85)
  );

  aliasv xaliasv84 (
	.PLUS(s_aib84),
	.MINUS(aib84)
  );

  aliasv xaliasv83 (
	.PLUS(s_aib83),
	.MINUS(aib83)
  );

  aliasv xaliasv82 (
	.PLUS(s_aib82),
	.MINUS(aib82)
  );

  aliasv xaliasv81 (
	.PLUS(s_aib81),
	.MINUS(aib81)
  );

  aliasv xaliasv80 (
	.PLUS(s_aib80),
	.MINUS(aib80)
  );

  aliasv xaliasv79 (
	.PLUS(s_aib79),
	.MINUS(aib79)
  );

  aliasv xaliasv78 (
	.PLUS(s_aib78),
	.MINUS(aib78)
  );

  aliasv xaliasv77 (
	.PLUS(s_aib77),
	.MINUS(aib77)
  );

  aliasv xaliasv76 (
	.PLUS(s_aib76),
	.MINUS(aib76)
  );

  aliasv xaliasv75 (
	.PLUS(s_aib75),
	.MINUS(aib75)
  );

  aliasv xaliasv74 (
	.PLUS(s_aib74),
	.MINUS(aib74)
  );

  aliasv xaliasv73 (
	.PLUS(s_aib73),
	.MINUS(aib73)
  );

  aliasv xaliasv72 (
	.PLUS(s_aib72),
	.MINUS(aib72)
  );

  aliasv xaliasv71 (
	.PLUS(s_aib71),
	.MINUS(aib71)
  );

  aliasv xaliasv70 (
	.PLUS(s_aib70),
	.MINUS(aib70)
  );

  aliasv xaliasv69 (
	.PLUS(s_aib69),
	.MINUS(aib69)
  );

  aliasv xaliasv68 (
	.PLUS(s_aib68),
	.MINUS(aib68)
  );

  aliasv xaliasv67 (
	.PLUS(s_aib67),
	.MINUS(aib67)
  );

  aliasv xaliasv66 (
	.PLUS(s_aib66),
	.MINUS(aib66)
  );

  aliasv xaliasv65 (
	.PLUS(s_aib65),
	.MINUS(aib65)
  );

  aliasv xaliasv64 (
	.PLUS(s_aib64),
	.MINUS(aib64)
  );

  aliasv xaliasv63 (
	.PLUS(s_aib63),
	.MINUS(aib63)
  );

  aliasv xaliasv62 (
	.PLUS(s_aib62),
	.MINUS(aib62)
  );

  aliasv xaliasv61 (
	.PLUS(s_aib61),
	.MINUS(aib61)
  );

  aliasv xaliasv60 (
	.PLUS(s_aib60),
	.MINUS(aib60)
  );

  aliasv xaliasv59 (
	.PLUS(s_aib59),
	.MINUS(aib59)
  );

  aliasv xaliasv58 (
	.PLUS(s_aib58),
	.MINUS(aib58)
  );

  aliasv xaliasv57 (
	.PLUS(s_aib57),
	.MINUS(aib57)
  );

  aliasv xaliasv56 (
	.PLUS(s_aib56),
	.MINUS(aib56)
  );

  aliasv xaliasv55 (
	.PLUS(s_aib55),
	.MINUS(aib55)
  );

  aliasv xaliasv54 (
	.PLUS(s_aib54),
	.MINUS(aib54)
  );

  aliasv xaliasv53 (
	.PLUS(s_aib53),
	.MINUS(aib53)
  );

  aliasv xaliasv52 (
	.PLUS(s_aib52),
	.MINUS(aib52)
  );

  aliasv xaliasv51 (
	.PLUS(s_aib51),
	.MINUS(aib51)
  );

  aliasv xaliasv50 (
	.PLUS(s_aib50),
	.MINUS(aib50)
  );

  aliasv xaliasv49 (
	.PLUS(s_aib49),
	.MINUS(aib49)
  );

  aliasv xaliasv48 (
	.PLUS(s_aib48),
	.MINUS(aib48)
  );

  aliasv xaliasv47 (
	.PLUS(s_aib47),
	.MINUS(aib47)
  );

  aliasv xaliasv46 (
	.PLUS(s_aib46),
	.MINUS(aib46)
  );

  aliasv xaliasv45 (
	.PLUS(s_aib45),
	.MINUS(aib45)
  );

  aliasv xaliasv44 (
	.PLUS(s_aib44),
	.MINUS(aib44)
  );

  aliasv xaliasv43 (
	.PLUS(s_aib43),
	.MINUS(aib43)
  );

  aliasv xaliasv42 (
	.PLUS(s_aib42),
	.MINUS(aib42)
  );

  aliasv xaliasv41 (
	.PLUS(s_aib41),
	.MINUS(aib41)
  );

  aliasv xaliasv40 (
	.PLUS(s_aib40),
	.MINUS(aib40)
  );

  aliasv xaliasv39 (
	.PLUS(s_aib39),
	.MINUS(aib39)
  );

  aliasv xaliasv38 (
	.PLUS(s_aib38),
	.MINUS(aib38)
  );

  aliasv xaliasv37 (
	.PLUS(s_aib37),
	.MINUS(aib37)
  );

  aliasv xaliasv36 (
	.PLUS(s_aib36),
	.MINUS(aib36)
  );

  aliasv xaliasv35 (
	.PLUS(s_aib35),
	.MINUS(aib35)
  );

  aliasv xaliasv34 (
	.PLUS(s_aib34),
	.MINUS(aib34)
  );

  aliasv xaliasv33 (
	.PLUS(s_aib33),
	.MINUS(aib33)
  );

  aliasv xaliasv32 (
	.PLUS(s_aib32),
	.MINUS(aib32)
  );

  aliasv xaliasv31 (
	.PLUS(s_aib31),
	.MINUS(aib31)
  );

  aliasv xaliasv30 (
	.PLUS(s_aib30),
	.MINUS(aib30)
  );

  aliasv xaliasv29 (
	.PLUS(s_aib29),
	.MINUS(aib29)
  );

  aliasv xaliasv28 (
	.PLUS(s_aib28),
	.MINUS(aib28)
  );

  aliasv xaliasv27 (
	.PLUS(s_aib27),
	.MINUS(aib27)
  );

  aliasv xaliasv26 (
	.PLUS(s_aib26),
	.MINUS(aib26)
  );

  aliasv xaliasv25 (
	.PLUS(s_aib25),
	.MINUS(aib25)
  );

  aliasv xaliasv24 (
	.PLUS(s_aib24),
	.MINUS(aib24)
  );

  aliasv xaliasv23 (
	.PLUS(s_aib23),
	.MINUS(aib23)
  );

  aliasv xaliasv22 (
	.PLUS(s_aib22),
	.MINUS(aib22)
  );

  aliasv xaliasv21 (
	.PLUS(s_aib21),
	.MINUS(aib21)
  );

  aliasv xaliasv20 (
	.PLUS(s_aib20),
	.MINUS(aib20)
  );

  aliasv xaliasv19 (
	.PLUS(s_aib19),
	.MINUS(aib19)
  );

  aliasv xaliasv18 (
	.PLUS(s_aib18),
	.MINUS(aib18)
  );

  aliasv xaliasv17 (
	.PLUS(s_aib17),
	.MINUS(aib17)
  );

  aliasv xaliasv16 (
	.PLUS(s_aib16),
	.MINUS(aib16)
  );

  aliasv xaliasv15 (
	.PLUS(s_aib15),
	.MINUS(aib15)
  );

  aliasv xaliasv14 (
	.PLUS(s_aib14),
	.MINUS(aib14)
  );

  aliasv xaliasv13 (
	.PLUS(s_aib13),
	.MINUS(aib13)
  );

  aliasv xaliasv12 (
	.PLUS(s_aib12),
	.MINUS(aib12)
  );

  aliasv xaliasv11 (
	.PLUS(s_aib11),
	.MINUS(aib11)
  );

  aliasv xaliasv10 (
	.PLUS(s_aib10),
	.MINUS(aib10)
  );

  aliasv xaliasv9 (
	.PLUS(s_aib9),
	.MINUS(aib9)
  );

  aliasv xaliasv8 (
	.PLUS(s_aib8),
	.MINUS(aib8)
  );

  aliasv xaliasv7 (
	.PLUS(s_aib7),
	.MINUS(aib7)
  );

  aliasv xaliasv6 (
	.PLUS(s_aib6),
	.MINUS(aib6)
  );

  aliasv xaliasv5 (
	.PLUS(s_aib5),
	.MINUS(aib5)
  );

  aliasv xaliasv4 (
	.PLUS(s_aib4),
	.MINUS(aib4)
  );

  aliasv xaliasv3 (
	.PLUS(s_aib3),
	.MINUS(aib3)
  );

  aliasv xaliasv2 (
	.PLUS(s_aib2),
	.MINUS(aib2)
  );

  aliasv xaliasv1 (
	.PLUS(s_aib1),
	.MINUS(aib1)
  );

  aliasv xaliasv0 (
	.PLUS(s_aib0),
	.MINUS(aib0)
  );


endmodule
