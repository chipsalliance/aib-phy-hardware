// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. 
// *****************************************************************************
// *****************************************************************************
//  Copyright © 2016 Altera Corporation. 
// *****************************************************************************
//  Module Name :  c3lib_ecc_dec_c88_d80
//  Date        :  Thu Jan 26 18:07:16 2017
//  Description :  ECC checker (based on the standard Extended Hamming Code
//                 scheme). Code generated by ecc_chk.pl script (command line
//                 options used: -num_data_bits 80).
// *****************************************************************************

module c3lib_ecc_dec_c88_d80(

  output logic		o_int_sec,
  output logic		o_int_ded,
  output logic[ 6 : 0 ]	o_syndrome,

  input  logic[ 87 : 0 ]	i_code,
  output logic[ 79 : 0 ]	o_data

);

// Declarations
var logic		parity0;
var logic[ 87 : 1 ]	correct_bit;

// Validate parity bits
assign parity0 = i_code[ 0 ] ^ i_code[ 1 ] ^ i_code[ 2 ] ^ i_code[ 3 ] ^ i_code[ 4 ] ^ i_code[ 5 ] ^ i_code[ 6 ] ^ i_code[ 7 ] ^ i_code[ 8 ] ^ i_code[ 9 ] ^ i_code[ 10 ] ^ i_code[ 11 ] ^ i_code[ 12 ] ^ i_code[ 13 ] ^ i_code[ 14 ] ^ i_code[ 15 ] ^ i_code[ 16 ] ^ i_code[ 17 ] ^ i_code[ 18 ] ^ i_code[ 19 ] ^ i_code[ 20 ] ^ i_code[ 21 ] ^ i_code[ 22 ] ^ i_code[ 23 ] ^ i_code[ 24 ] ^ i_code[ 25 ] ^ i_code[ 26 ] ^ i_code[ 27 ] ^ i_code[ 28 ] ^ i_code[ 29 ] ^ i_code[ 30 ] ^ i_code[ 31 ] ^ i_code[ 32 ] ^ i_code[ 33 ] ^ i_code[ 34 ] ^ i_code[ 35 ] ^ i_code[ 36 ] ^ i_code[ 37 ] ^ i_code[ 38 ] ^ i_code[ 39 ] ^ i_code[ 40 ] ^ i_code[ 41 ] ^ i_code[ 42 ] ^ i_code[ 43 ] ^ i_code[ 44 ] ^ i_code[ 45 ] ^ i_code[ 46 ] ^ i_code[ 47 ] ^ i_code[ 48 ] ^ i_code[ 49 ] ^ i_code[ 50 ] ^ i_code[ 51 ] ^ i_code[ 52 ] ^ i_code[ 53 ] ^ i_code[ 54 ] ^ i_code[ 55 ] ^ i_code[ 56 ] ^ i_code[ 57 ] ^ i_code[ 58 ] ^ i_code[ 59 ] ^ i_code[ 60 ] ^ i_code[ 61 ] ^ i_code[ 62 ] ^ i_code[ 63 ] ^ i_code[ 64 ] ^ i_code[ 65 ] ^ i_code[ 66 ] ^ i_code[ 67 ] ^ i_code[ 68 ] ^ i_code[ 69 ] ^ i_code[ 70 ] ^ i_code[ 71 ] ^ i_code[ 72 ] ^ i_code[ 73 ] ^ i_code[ 74 ] ^ i_code[ 75 ] ^ i_code[ 76 ] ^ i_code[ 77 ] ^ i_code[ 78 ] ^ i_code[ 79 ] ^ i_code[ 80 ] ^ i_code[ 81 ] ^ i_code[ 82 ] ^ i_code[ 83 ] ^ i_code[ 84 ] ^ i_code[ 85 ] ^ i_code[ 86 ] ^ i_code[ 87 ];
assign o_syndrome[ 0 ] = i_code[ 1 ] ^ i_code[ 3 ] ^ i_code[ 5 ] ^ i_code[ 7 ] ^ i_code[ 9 ] ^ i_code[ 11 ] ^ i_code[ 13 ] ^ i_code[ 15 ] ^ i_code[ 17 ] ^ i_code[ 19 ] ^ i_code[ 21 ] ^ i_code[ 23 ] ^ i_code[ 25 ] ^ i_code[ 27 ] ^ i_code[ 29 ] ^ i_code[ 31 ] ^ i_code[ 33 ] ^ i_code[ 35 ] ^ i_code[ 37 ] ^ i_code[ 39 ] ^ i_code[ 41 ] ^ i_code[ 43 ] ^ i_code[ 45 ] ^ i_code[ 47 ] ^ i_code[ 49 ] ^ i_code[ 51 ] ^ i_code[ 53 ] ^ i_code[ 55 ] ^ i_code[ 57 ] ^ i_code[ 59 ] ^ i_code[ 61 ] ^ i_code[ 63 ] ^ i_code[ 65 ] ^ i_code[ 67 ] ^ i_code[ 69 ] ^ i_code[ 71 ] ^ i_code[ 73 ] ^ i_code[ 75 ] ^ i_code[ 77 ] ^ i_code[ 79 ] ^ i_code[ 81 ] ^ i_code[ 83 ] ^ i_code[ 85 ] ^ i_code[ 87 ];
assign o_syndrome[ 1 ] = i_code[ 2 ] ^ i_code[ 3 ] ^ i_code[ 6 ] ^ i_code[ 7 ] ^ i_code[ 10 ] ^ i_code[ 11 ] ^ i_code[ 14 ] ^ i_code[ 15 ] ^ i_code[ 18 ] ^ i_code[ 19 ] ^ i_code[ 22 ] ^ i_code[ 23 ] ^ i_code[ 26 ] ^ i_code[ 27 ] ^ i_code[ 30 ] ^ i_code[ 31 ] ^ i_code[ 34 ] ^ i_code[ 35 ] ^ i_code[ 38 ] ^ i_code[ 39 ] ^ i_code[ 42 ] ^ i_code[ 43 ] ^ i_code[ 46 ] ^ i_code[ 47 ] ^ i_code[ 50 ] ^ i_code[ 51 ] ^ i_code[ 54 ] ^ i_code[ 55 ] ^ i_code[ 58 ] ^ i_code[ 59 ] ^ i_code[ 62 ] ^ i_code[ 63 ] ^ i_code[ 66 ] ^ i_code[ 67 ] ^ i_code[ 70 ] ^ i_code[ 71 ] ^ i_code[ 74 ] ^ i_code[ 75 ] ^ i_code[ 78 ] ^ i_code[ 79 ] ^ i_code[ 82 ] ^ i_code[ 83 ] ^ i_code[ 86 ] ^ i_code[ 87 ];
assign o_syndrome[ 2 ] = i_code[ 4 ] ^ i_code[ 5 ] ^ i_code[ 6 ] ^ i_code[ 7 ] ^ i_code[ 12 ] ^ i_code[ 13 ] ^ i_code[ 14 ] ^ i_code[ 15 ] ^ i_code[ 20 ] ^ i_code[ 21 ] ^ i_code[ 22 ] ^ i_code[ 23 ] ^ i_code[ 28 ] ^ i_code[ 29 ] ^ i_code[ 30 ] ^ i_code[ 31 ] ^ i_code[ 36 ] ^ i_code[ 37 ] ^ i_code[ 38 ] ^ i_code[ 39 ] ^ i_code[ 44 ] ^ i_code[ 45 ] ^ i_code[ 46 ] ^ i_code[ 47 ] ^ i_code[ 52 ] ^ i_code[ 53 ] ^ i_code[ 54 ] ^ i_code[ 55 ] ^ i_code[ 60 ] ^ i_code[ 61 ] ^ i_code[ 62 ] ^ i_code[ 63 ] ^ i_code[ 68 ] ^ i_code[ 69 ] ^ i_code[ 70 ] ^ i_code[ 71 ] ^ i_code[ 76 ] ^ i_code[ 77 ] ^ i_code[ 78 ] ^ i_code[ 79 ] ^ i_code[ 84 ] ^ i_code[ 85 ] ^ i_code[ 86 ] ^ i_code[ 87 ];
assign o_syndrome[ 3 ] = i_code[ 8 ] ^ i_code[ 9 ] ^ i_code[ 10 ] ^ i_code[ 11 ] ^ i_code[ 12 ] ^ i_code[ 13 ] ^ i_code[ 14 ] ^ i_code[ 15 ] ^ i_code[ 24 ] ^ i_code[ 25 ] ^ i_code[ 26 ] ^ i_code[ 27 ] ^ i_code[ 28 ] ^ i_code[ 29 ] ^ i_code[ 30 ] ^ i_code[ 31 ] ^ i_code[ 40 ] ^ i_code[ 41 ] ^ i_code[ 42 ] ^ i_code[ 43 ] ^ i_code[ 44 ] ^ i_code[ 45 ] ^ i_code[ 46 ] ^ i_code[ 47 ] ^ i_code[ 56 ] ^ i_code[ 57 ] ^ i_code[ 58 ] ^ i_code[ 59 ] ^ i_code[ 60 ] ^ i_code[ 61 ] ^ i_code[ 62 ] ^ i_code[ 63 ] ^ i_code[ 72 ] ^ i_code[ 73 ] ^ i_code[ 74 ] ^ i_code[ 75 ] ^ i_code[ 76 ] ^ i_code[ 77 ] ^ i_code[ 78 ] ^ i_code[ 79 ];
assign o_syndrome[ 4 ] = i_code[ 16 ] ^ i_code[ 17 ] ^ i_code[ 18 ] ^ i_code[ 19 ] ^ i_code[ 20 ] ^ i_code[ 21 ] ^ i_code[ 22 ] ^ i_code[ 23 ] ^ i_code[ 24 ] ^ i_code[ 25 ] ^ i_code[ 26 ] ^ i_code[ 27 ] ^ i_code[ 28 ] ^ i_code[ 29 ] ^ i_code[ 30 ] ^ i_code[ 31 ] ^ i_code[ 48 ] ^ i_code[ 49 ] ^ i_code[ 50 ] ^ i_code[ 51 ] ^ i_code[ 52 ] ^ i_code[ 53 ] ^ i_code[ 54 ] ^ i_code[ 55 ] ^ i_code[ 56 ] ^ i_code[ 57 ] ^ i_code[ 58 ] ^ i_code[ 59 ] ^ i_code[ 60 ] ^ i_code[ 61 ] ^ i_code[ 62 ] ^ i_code[ 63 ] ^ i_code[ 80 ] ^ i_code[ 81 ] ^ i_code[ 82 ] ^ i_code[ 83 ] ^ i_code[ 84 ] ^ i_code[ 85 ] ^ i_code[ 86 ] ^ i_code[ 87 ];
assign o_syndrome[ 5 ] = i_code[ 32 ] ^ i_code[ 33 ] ^ i_code[ 34 ] ^ i_code[ 35 ] ^ i_code[ 36 ] ^ i_code[ 37 ] ^ i_code[ 38 ] ^ i_code[ 39 ] ^ i_code[ 40 ] ^ i_code[ 41 ] ^ i_code[ 42 ] ^ i_code[ 43 ] ^ i_code[ 44 ] ^ i_code[ 45 ] ^ i_code[ 46 ] ^ i_code[ 47 ] ^ i_code[ 48 ] ^ i_code[ 49 ] ^ i_code[ 50 ] ^ i_code[ 51 ] ^ i_code[ 52 ] ^ i_code[ 53 ] ^ i_code[ 54 ] ^ i_code[ 55 ] ^ i_code[ 56 ] ^ i_code[ 57 ] ^ i_code[ 58 ] ^ i_code[ 59 ] ^ i_code[ 60 ] ^ i_code[ 61 ] ^ i_code[ 62 ] ^ i_code[ 63 ];
assign o_syndrome[ 6 ] = i_code[ 64 ] ^ i_code[ 65 ] ^ i_code[ 66 ] ^ i_code[ 67 ] ^ i_code[ 68 ] ^ i_code[ 69 ] ^ i_code[ 70 ] ^ i_code[ 71 ] ^ i_code[ 72 ] ^ i_code[ 73 ] ^ i_code[ 74 ] ^ i_code[ 75 ] ^ i_code[ 76 ] ^ i_code[ 77 ] ^ i_code[ 78 ] ^ i_code[ 79 ] ^ i_code[ 80 ] ^ i_code[ 81 ] ^ i_code[ 82 ] ^ i_code[ 83 ] ^ i_code[ 84 ] ^ i_code[ 85 ] ^ i_code[ 86 ] ^ i_code[ 87 ];

// Decision logic
assign o_int_sec  = parity0;
assign o_int_ded  = !parity0 && (|o_syndrome);
assign correct_bit[ 1 ] = (o_syndrome == 7'd1);
assign correct_bit[ 2 ] = (o_syndrome == 7'd2);
assign correct_bit[ 3 ] = (o_syndrome == 7'd3);
assign correct_bit[ 4 ] = (o_syndrome == 7'd4);
assign correct_bit[ 5 ] = (o_syndrome == 7'd5);
assign correct_bit[ 6 ] = (o_syndrome == 7'd6);
assign correct_bit[ 7 ] = (o_syndrome == 7'd7);
assign correct_bit[ 8 ] = (o_syndrome == 7'd8);
assign correct_bit[ 9 ] = (o_syndrome == 7'd9);
assign correct_bit[ 10 ] = (o_syndrome == 7'd10);
assign correct_bit[ 11 ] = (o_syndrome == 7'd11);
assign correct_bit[ 12 ] = (o_syndrome == 7'd12);
assign correct_bit[ 13 ] = (o_syndrome == 7'd13);
assign correct_bit[ 14 ] = (o_syndrome == 7'd14);
assign correct_bit[ 15 ] = (o_syndrome == 7'd15);
assign correct_bit[ 16 ] = (o_syndrome == 7'd16);
assign correct_bit[ 17 ] = (o_syndrome == 7'd17);
assign correct_bit[ 18 ] = (o_syndrome == 7'd18);
assign correct_bit[ 19 ] = (o_syndrome == 7'd19);
assign correct_bit[ 20 ] = (o_syndrome == 7'd20);
assign correct_bit[ 21 ] = (o_syndrome == 7'd21);
assign correct_bit[ 22 ] = (o_syndrome == 7'd22);
assign correct_bit[ 23 ] = (o_syndrome == 7'd23);
assign correct_bit[ 24 ] = (o_syndrome == 7'd24);
assign correct_bit[ 25 ] = (o_syndrome == 7'd25);
assign correct_bit[ 26 ] = (o_syndrome == 7'd26);
assign correct_bit[ 27 ] = (o_syndrome == 7'd27);
assign correct_bit[ 28 ] = (o_syndrome == 7'd28);
assign correct_bit[ 29 ] = (o_syndrome == 7'd29);
assign correct_bit[ 30 ] = (o_syndrome == 7'd30);
assign correct_bit[ 31 ] = (o_syndrome == 7'd31);
assign correct_bit[ 32 ] = (o_syndrome == 7'd32);
assign correct_bit[ 33 ] = (o_syndrome == 7'd33);
assign correct_bit[ 34 ] = (o_syndrome == 7'd34);
assign correct_bit[ 35 ] = (o_syndrome == 7'd35);
assign correct_bit[ 36 ] = (o_syndrome == 7'd36);
assign correct_bit[ 37 ] = (o_syndrome == 7'd37);
assign correct_bit[ 38 ] = (o_syndrome == 7'd38);
assign correct_bit[ 39 ] = (o_syndrome == 7'd39);
assign correct_bit[ 40 ] = (o_syndrome == 7'd40);
assign correct_bit[ 41 ] = (o_syndrome == 7'd41);
assign correct_bit[ 42 ] = (o_syndrome == 7'd42);
assign correct_bit[ 43 ] = (o_syndrome == 7'd43);
assign correct_bit[ 44 ] = (o_syndrome == 7'd44);
assign correct_bit[ 45 ] = (o_syndrome == 7'd45);
assign correct_bit[ 46 ] = (o_syndrome == 7'd46);
assign correct_bit[ 47 ] = (o_syndrome == 7'd47);
assign correct_bit[ 48 ] = (o_syndrome == 7'd48);
assign correct_bit[ 49 ] = (o_syndrome == 7'd49);
assign correct_bit[ 50 ] = (o_syndrome == 7'd50);
assign correct_bit[ 51 ] = (o_syndrome == 7'd51);
assign correct_bit[ 52 ] = (o_syndrome == 7'd52);
assign correct_bit[ 53 ] = (o_syndrome == 7'd53);
assign correct_bit[ 54 ] = (o_syndrome == 7'd54);
assign correct_bit[ 55 ] = (o_syndrome == 7'd55);
assign correct_bit[ 56 ] = (o_syndrome == 7'd56);
assign correct_bit[ 57 ] = (o_syndrome == 7'd57);
assign correct_bit[ 58 ] = (o_syndrome == 7'd58);
assign correct_bit[ 59 ] = (o_syndrome == 7'd59);
assign correct_bit[ 60 ] = (o_syndrome == 7'd60);
assign correct_bit[ 61 ] = (o_syndrome == 7'd61);
assign correct_bit[ 62 ] = (o_syndrome == 7'd62);
assign correct_bit[ 63 ] = (o_syndrome == 7'd63);
assign correct_bit[ 64 ] = (o_syndrome == 7'd64);
assign correct_bit[ 65 ] = (o_syndrome == 7'd65);
assign correct_bit[ 66 ] = (o_syndrome == 7'd66);
assign correct_bit[ 67 ] = (o_syndrome == 7'd67);
assign correct_bit[ 68 ] = (o_syndrome == 7'd68);
assign correct_bit[ 69 ] = (o_syndrome == 7'd69);
assign correct_bit[ 70 ] = (o_syndrome == 7'd70);
assign correct_bit[ 71 ] = (o_syndrome == 7'd71);
assign correct_bit[ 72 ] = (o_syndrome == 7'd72);
assign correct_bit[ 73 ] = (o_syndrome == 7'd73);
assign correct_bit[ 74 ] = (o_syndrome == 7'd74);
assign correct_bit[ 75 ] = (o_syndrome == 7'd75);
assign correct_bit[ 76 ] = (o_syndrome == 7'd76);
assign correct_bit[ 77 ] = (o_syndrome == 7'd77);
assign correct_bit[ 78 ] = (o_syndrome == 7'd78);
assign correct_bit[ 79 ] = (o_syndrome == 7'd79);
assign correct_bit[ 80 ] = (o_syndrome == 7'd80);
assign correct_bit[ 81 ] = (o_syndrome == 7'd81);
assign correct_bit[ 82 ] = (o_syndrome == 7'd82);
assign correct_bit[ 83 ] = (o_syndrome == 7'd83);
assign correct_bit[ 84 ] = (o_syndrome == 7'd84);
assign correct_bit[ 85 ] = (o_syndrome == 7'd85);
assign correct_bit[ 86 ] = (o_syndrome == 7'd86);
assign correct_bit[ 87 ] = (o_syndrome == 7'd87);

// Extract data bits
assign o_data[ 0 ] = correct_bit[ 3 ]? ~i_code[ 3 ] : i_code[ 3 ];
assign o_data[ 1 ] = correct_bit[ 5 ]? ~i_code[ 5 ] : i_code[ 5 ];
assign o_data[ 2 ] = correct_bit[ 6 ]? ~i_code[ 6 ] : i_code[ 6 ];
assign o_data[ 3 ] = correct_bit[ 7 ]? ~i_code[ 7 ] : i_code[ 7 ];
assign o_data[ 4 ] = correct_bit[ 9 ]? ~i_code[ 9 ] : i_code[ 9 ];
assign o_data[ 5 ] = correct_bit[ 10 ]? ~i_code[ 10 ] : i_code[ 10 ];
assign o_data[ 6 ] = correct_bit[ 11 ]? ~i_code[ 11 ] : i_code[ 11 ];
assign o_data[ 7 ] = correct_bit[ 12 ]? ~i_code[ 12 ] : i_code[ 12 ];
assign o_data[ 8 ] = correct_bit[ 13 ]? ~i_code[ 13 ] : i_code[ 13 ];
assign o_data[ 9 ] = correct_bit[ 14 ]? ~i_code[ 14 ] : i_code[ 14 ];
assign o_data[ 10 ] = correct_bit[ 15 ]? ~i_code[ 15 ] : i_code[ 15 ];
assign o_data[ 11 ] = correct_bit[ 17 ]? ~i_code[ 17 ] : i_code[ 17 ];
assign o_data[ 12 ] = correct_bit[ 18 ]? ~i_code[ 18 ] : i_code[ 18 ];
assign o_data[ 13 ] = correct_bit[ 19 ]? ~i_code[ 19 ] : i_code[ 19 ];
assign o_data[ 14 ] = correct_bit[ 20 ]? ~i_code[ 20 ] : i_code[ 20 ];
assign o_data[ 15 ] = correct_bit[ 21 ]? ~i_code[ 21 ] : i_code[ 21 ];
assign o_data[ 16 ] = correct_bit[ 22 ]? ~i_code[ 22 ] : i_code[ 22 ];
assign o_data[ 17 ] = correct_bit[ 23 ]? ~i_code[ 23 ] : i_code[ 23 ];
assign o_data[ 18 ] = correct_bit[ 24 ]? ~i_code[ 24 ] : i_code[ 24 ];
assign o_data[ 19 ] = correct_bit[ 25 ]? ~i_code[ 25 ] : i_code[ 25 ];
assign o_data[ 20 ] = correct_bit[ 26 ]? ~i_code[ 26 ] : i_code[ 26 ];
assign o_data[ 21 ] = correct_bit[ 27 ]? ~i_code[ 27 ] : i_code[ 27 ];
assign o_data[ 22 ] = correct_bit[ 28 ]? ~i_code[ 28 ] : i_code[ 28 ];
assign o_data[ 23 ] = correct_bit[ 29 ]? ~i_code[ 29 ] : i_code[ 29 ];
assign o_data[ 24 ] = correct_bit[ 30 ]? ~i_code[ 30 ] : i_code[ 30 ];
assign o_data[ 25 ] = correct_bit[ 31 ]? ~i_code[ 31 ] : i_code[ 31 ];
assign o_data[ 26 ] = correct_bit[ 33 ]? ~i_code[ 33 ] : i_code[ 33 ];
assign o_data[ 27 ] = correct_bit[ 34 ]? ~i_code[ 34 ] : i_code[ 34 ];
assign o_data[ 28 ] = correct_bit[ 35 ]? ~i_code[ 35 ] : i_code[ 35 ];
assign o_data[ 29 ] = correct_bit[ 36 ]? ~i_code[ 36 ] : i_code[ 36 ];
assign o_data[ 30 ] = correct_bit[ 37 ]? ~i_code[ 37 ] : i_code[ 37 ];
assign o_data[ 31 ] = correct_bit[ 38 ]? ~i_code[ 38 ] : i_code[ 38 ];
assign o_data[ 32 ] = correct_bit[ 39 ]? ~i_code[ 39 ] : i_code[ 39 ];
assign o_data[ 33 ] = correct_bit[ 40 ]? ~i_code[ 40 ] : i_code[ 40 ];
assign o_data[ 34 ] = correct_bit[ 41 ]? ~i_code[ 41 ] : i_code[ 41 ];
assign o_data[ 35 ] = correct_bit[ 42 ]? ~i_code[ 42 ] : i_code[ 42 ];
assign o_data[ 36 ] = correct_bit[ 43 ]? ~i_code[ 43 ] : i_code[ 43 ];
assign o_data[ 37 ] = correct_bit[ 44 ]? ~i_code[ 44 ] : i_code[ 44 ];
assign o_data[ 38 ] = correct_bit[ 45 ]? ~i_code[ 45 ] : i_code[ 45 ];
assign o_data[ 39 ] = correct_bit[ 46 ]? ~i_code[ 46 ] : i_code[ 46 ];
assign o_data[ 40 ] = correct_bit[ 47 ]? ~i_code[ 47 ] : i_code[ 47 ];
assign o_data[ 41 ] = correct_bit[ 48 ]? ~i_code[ 48 ] : i_code[ 48 ];
assign o_data[ 42 ] = correct_bit[ 49 ]? ~i_code[ 49 ] : i_code[ 49 ];
assign o_data[ 43 ] = correct_bit[ 50 ]? ~i_code[ 50 ] : i_code[ 50 ];
assign o_data[ 44 ] = correct_bit[ 51 ]? ~i_code[ 51 ] : i_code[ 51 ];
assign o_data[ 45 ] = correct_bit[ 52 ]? ~i_code[ 52 ] : i_code[ 52 ];
assign o_data[ 46 ] = correct_bit[ 53 ]? ~i_code[ 53 ] : i_code[ 53 ];
assign o_data[ 47 ] = correct_bit[ 54 ]? ~i_code[ 54 ] : i_code[ 54 ];
assign o_data[ 48 ] = correct_bit[ 55 ]? ~i_code[ 55 ] : i_code[ 55 ];
assign o_data[ 49 ] = correct_bit[ 56 ]? ~i_code[ 56 ] : i_code[ 56 ];
assign o_data[ 50 ] = correct_bit[ 57 ]? ~i_code[ 57 ] : i_code[ 57 ];
assign o_data[ 51 ] = correct_bit[ 58 ]? ~i_code[ 58 ] : i_code[ 58 ];
assign o_data[ 52 ] = correct_bit[ 59 ]? ~i_code[ 59 ] : i_code[ 59 ];
assign o_data[ 53 ] = correct_bit[ 60 ]? ~i_code[ 60 ] : i_code[ 60 ];
assign o_data[ 54 ] = correct_bit[ 61 ]? ~i_code[ 61 ] : i_code[ 61 ];
assign o_data[ 55 ] = correct_bit[ 62 ]? ~i_code[ 62 ] : i_code[ 62 ];
assign o_data[ 56 ] = correct_bit[ 63 ]? ~i_code[ 63 ] : i_code[ 63 ];
assign o_data[ 57 ] = correct_bit[ 65 ]? ~i_code[ 65 ] : i_code[ 65 ];
assign o_data[ 58 ] = correct_bit[ 66 ]? ~i_code[ 66 ] : i_code[ 66 ];
assign o_data[ 59 ] = correct_bit[ 67 ]? ~i_code[ 67 ] : i_code[ 67 ];
assign o_data[ 60 ] = correct_bit[ 68 ]? ~i_code[ 68 ] : i_code[ 68 ];
assign o_data[ 61 ] = correct_bit[ 69 ]? ~i_code[ 69 ] : i_code[ 69 ];
assign o_data[ 62 ] = correct_bit[ 70 ]? ~i_code[ 70 ] : i_code[ 70 ];
assign o_data[ 63 ] = correct_bit[ 71 ]? ~i_code[ 71 ] : i_code[ 71 ];
assign o_data[ 64 ] = correct_bit[ 72 ]? ~i_code[ 72 ] : i_code[ 72 ];
assign o_data[ 65 ] = correct_bit[ 73 ]? ~i_code[ 73 ] : i_code[ 73 ];
assign o_data[ 66 ] = correct_bit[ 74 ]? ~i_code[ 74 ] : i_code[ 74 ];
assign o_data[ 67 ] = correct_bit[ 75 ]? ~i_code[ 75 ] : i_code[ 75 ];
assign o_data[ 68 ] = correct_bit[ 76 ]? ~i_code[ 76 ] : i_code[ 76 ];
assign o_data[ 69 ] = correct_bit[ 77 ]? ~i_code[ 77 ] : i_code[ 77 ];
assign o_data[ 70 ] = correct_bit[ 78 ]? ~i_code[ 78 ] : i_code[ 78 ];
assign o_data[ 71 ] = correct_bit[ 79 ]? ~i_code[ 79 ] : i_code[ 79 ];
assign o_data[ 72 ] = correct_bit[ 80 ]? ~i_code[ 80 ] : i_code[ 80 ];
assign o_data[ 73 ] = correct_bit[ 81 ]? ~i_code[ 81 ] : i_code[ 81 ];
assign o_data[ 74 ] = correct_bit[ 82 ]? ~i_code[ 82 ] : i_code[ 82 ];
assign o_data[ 75 ] = correct_bit[ 83 ]? ~i_code[ 83 ] : i_code[ 83 ];
assign o_data[ 76 ] = correct_bit[ 84 ]? ~i_code[ 84 ] : i_code[ 84 ];
assign o_data[ 77 ] = correct_bit[ 85 ]? ~i_code[ 85 ] : i_code[ 85 ];
assign o_data[ 78 ] = correct_bit[ 86 ]? ~i_code[ 86 ] : i_code[ 86 ];
assign o_data[ 79 ] = correct_bit[ 87 ]? ~i_code[ 87 ] : i_code[ 87 ];

endmodule

