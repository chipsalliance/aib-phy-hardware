// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. All rights reserved
module aibcr3_aliasd(ra, rb);
 input ra;
 output rb;
  assign rb = ra;
endmodule




