// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. All rights reserved


module aibnd_fine_dly_x1 ( sp,sn , dout); // vcc_regphy, vss_io );

  input sp,sn;
  output dout;
//  input vss_io;
//  input vcc_regphy;


  assign dout = 1'bz ;

endmodule


