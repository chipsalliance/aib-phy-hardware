// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. 
// Library - aibnd_lib, Cell - aibnd_d8xsesdd2, View - schematic
// LAST TIME SAVED: Nov 20 19:10:52 2014
// NETLIST TIME: Nov 21 11:04:30 2014

module aibnd_d8xsesdd2 ( iopad, vccl_aibnd, vssl_aibnd );

inout  iopad;

input  vccl_aibnd, vssl_aibnd;

/*
specify 
    specparam CDS_LIBNAME  = "aibnd_lib";
    specparam CDS_CELLNAME = "aibnd_d8xsesdd2";
    specparam CDS_VIEWNAME = "schematic";
endspecify
*/



endmodule

