// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. 
//------------------------------------------------------------------------
// Copyright (c) 2012 Altera Corporation. .
// Library - aibndaux_lib, Cell - aibndaux_async, View - schematic
// LAST TIME SAVED: Jul  8 16:37:33 2015
// NETLIST TIME: Jul  9 10:28:17 2015
// `timescale 1ns / 1ns 

module aibndaux_async ( io_out, jtag_rx_scan_out_10x7,
     jtag_rx_scan_out_10x8, last_bs_out_10x7, last_bs_out_10x8, tstmx,
     iopad_auxactred1, iopad_auxactred2, iopad_io_in, iopad_io_oe,
     iopad_io_out, iopad_tstmx, anlg_rstb, csr_actreden,
     csr_asyn_dataselb, csr_asyn_ndrv, csr_asyn_pdrv, csr_asyn_rxen,
     csr_asyn_txen, csr_iocsr_sel, dig_rstb, io_in, io_oe,
     jtag_clkdr_in5l, jtag_clkdr_in5r, jtag_clkdr_in6l,
     jtag_clkdr_in6r, jtag_clkdr_in7r, jtag_clkdr_in8r, jtag_clksel,
     jtag_intest, jtag_mode_in, jtag_rstb, jtag_rstb_en,
     jtag_tx_scan_in_01x5, jtag_tx_scan_in_01x6, jtag_tx_scanen_in,
     jtag_weakpdn, jtag_weakpu, last_bs_in_01x5, last_bs_in_01x6,
     crete_detect, vccl_aibndaux, vssl_aibndaux );

output  jtag_rx_scan_out_10x7, jtag_rx_scan_out_10x8, last_bs_out_10x7,
     last_bs_out_10x8;

inout  iopad_auxactred1, iopad_auxactred2;

input  anlg_rstb, csr_asyn_dataselb, csr_asyn_txen, csr_iocsr_sel,
     dig_rstb, jtag_clkdr_in5l, jtag_clkdr_in5r, jtag_clkdr_in6l,
     jtag_clkdr_in6r, jtag_clkdr_in7r, jtag_clkdr_in8r, jtag_clksel,
     jtag_intest, jtag_mode_in, jtag_rstb, jtag_rstb_en,
     jtag_tx_scan_in_01x5, jtag_tx_scan_in_01x6, jtag_tx_scanen_in,
     jtag_weakpdn, jtag_weakpu, last_bs_in_01x5, last_bs_in_01x6,
     crete_detect, vccl_aibndaux, vssl_aibndaux;

output [7:0]  tstmx;
output [7:0]  io_out;

inout [1:0]  iopad_io_oe;
inout [7:0]  iopad_tstmx;
inout [7:0]  iopad_io_out;
inout [7:0]  iopad_io_in;

input [2:0]  csr_asyn_rxen;
input [1:0]  csr_asyn_ndrv;
input [1:0]  io_oe;
input [12:0]  csr_actreden;
input [7:0]  io_in;
input [1:0]  csr_asyn_pdrv;

wire csr_iocsr_sel; // Conversion Sript Generated

// Buses in the design

wire  [2:0]  csr_asyn_rxen_int;

wire  [1:0]  csr_asyn_ndrv_int;

wire  [1:0]  csr_asyn_pdrv_int;


// specify 
//     specparam CDS_LIBNAME  = "aibndaux_lib";
//     specparam CDS_CELLNAME = "aibndaux_async";
//     specparam CDS_VIEWNAME = "schematic";
// endspecify

aibnd_buffx1_top  xauxactred1 ( .idata1_in1_jtag_out(net0624),
     .async_dat_in1_jtag_out(net0625), .idata0_in1_jtag_out(net0758),
     .prev_io_shift_en(csr_actreden[12]), .jtag_clkdr_outn(net0511),
     .anlg_rstb(anlg_rstb), .pd_data_aib(net0646), .oclk_out(net0633),
     .oclkb_out(net0606), .odat0_out(net0677), .odat1_out(net0647),
     .odat_async_out(auxactred1), .pd_data_out(net0700),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0({vssl_aibndaux, vccl_aibndaux, vssl_aibndaux}),
     .irxen_in1(csr_asyn_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(auxactred1_to_tstmx6), .oclkb_in1(vssl_aibndaux),
     .jtag_clksel(jtag_clksel), .odat0_in1(vssl_aibndaux),
     .vssl_aibnd(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(csr_actreden[12]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0601), .jtag_intest(jtag_intest),
     .odat1_aib(net0699), .jtag_rx_scan_out(jtag_rx_scan_out_10x8),
     .odat0_aib(net0675), .oclk_aib(net0701),
     .last_bs_out(last_bs_out_10x8), .vccl_aibnd(vccl_aibndaux),
     .oclkb_aib(net0693), .jtag_clkdr_in(jtag_clkdr_in8r),
     .jtag_rstb_en(jtag_rstb_en), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_in_11x8),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_11x8), .iopad(iopad_auxactred1),
     .oclkn(net0602), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xauxactred2 ( .idata1_in1_jtag_out(net0630),
     .async_dat_in1_jtag_out(net0631), .idata0_in1_jtag_out(net0748),
     .prev_io_shift_en(csr_actreden[12]), .jtag_clkdr_outn(net0512),
     .anlg_rstb(anlg_rstb), .pd_data_aib(net0626), .oclk_out(net0614),
     .oclkb_out(net0680), .odat0_out(net0702), .odat1_out(net0619),
     .odat_async_out(auxactred2), .pd_data_out(net0650),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0({vssl_aibndaux, vccl_aibndaux, vssl_aibndaux}),
     .irxen_in1(csr_asyn_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(auxactred2_to_tstmx7), .oclkb_in1(vssl_aibndaux),
     .jtag_clksel(jtag_clksel), .odat0_in1(vssl_aibndaux),
     .vssl_aibnd(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(csr_actreden[12]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0622), .jtag_intest(jtag_intest),
     .odat1_aib(net0692), .jtag_rx_scan_out(jtag_rx_scan_out_10x7),
     .odat0_aib(net0683), .oclk_aib(net0698),
     .last_bs_out(last_bs_out_10x7), .vccl_aibnd(vccl_aibndaux),
     .oclkb_aib(net0661), .jtag_clkdr_in(jtag_clkdr_in7r),
     .jtag_rstb_en(jtag_rstb_en), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_in_11x7),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_11x7), .iopad(iopad_auxactred2),
     .oclkn(net0629), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xtstmx4 ( .idata1_in1_jtag_out(net0744),
     .async_dat_in1_jtag_out(net0818), .idata0_in1_jtag_out(net0708),
     .prev_io_shift_en(csr_actreden[10]), .jtag_clkdr_outn(net0513),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(jtag_intest), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(jtag_rstb_en), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0663), .oclk_out(net0639), .oclkb_out(net0671),
     .odat0_out(net0649), .odat1_out(net0656),
     .odat_async_out(tstmx[4]), .pd_data_out(net0672),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0(csr_asyn_rxen_int[2:0]),
     .irxen_in1(csr_asyn_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(tstmx4_to_tstmx2), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(tstmx6_to_tstmx4), .shift_en(csr_actreden[11]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0160), .odat1_aib(net0673),
     .jtag_rx_scan_out(jtag_rx_scan_in_12x8), .odat0_aib(net0654),
     .oclk_aib(net0664), .last_bs_out(last_bs_in_12x8),
     .oclkb_aib(net0670), .jtag_clkdr_in(jtag_clkdr_in6r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_12x6),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_12x6), .iopad(iopad_tstmx[4]),
     .oclkn(net0660), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xtstmx5 ( .idata1_in1_jtag_out(net0718),
     .async_dat_in1_jtag_out(net0713), .idata0_in1_jtag_out(net0773),
     .prev_io_shift_en(csr_actreden[10]), .jtag_clkdr_outn(net0514),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(jtag_intest), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(jtag_rstb_en), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0645), .oclk_out(net0674), .oclkb_out(net0637),
     .odat0_out(net0644), .odat1_out(net0651),
     .odat_async_out(tstmx[5]), .pd_data_out(net0667),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0(csr_asyn_rxen_int[2:0]),
     .irxen_in1(csr_asyn_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(tstmx5_to_tstmx3), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(tstmx7_to_tstmx5), .shift_en(csr_actreden[11]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0153), .odat1_aib(net0669),
     .jtag_rx_scan_out(jtag_rx_scan_in_12x7), .odat0_aib(net0643),
     .oclk_aib(net0635), .last_bs_out(last_bs_in_12x7),
     .oclkb_aib(net0668), .jtag_clkdr_in(jtag_clkdr_in5r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_12x5),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_12x5), .iopad(iopad_tstmx[5]),
     .oclkn(net0665), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xtstmx2 ( .idata1_in1_jtag_out(net0722),
     .async_dat_in1_jtag_out(net0222), .idata0_in1_jtag_out(net0811),
     .prev_io_shift_en(csr_actreden[9]), .jtag_clkdr_outn(net0515),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(jtag_intest), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(jtag_rstb_en), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0342), .oclk_out(net0652), .oclkb_out(net0332),
     .odat0_out(net0333), .odat1_out(net0334),
     .odat_async_out(tstmx[2]), .pd_data_out(net0335),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0(csr_asyn_rxen_int[2:0]),
     .irxen_in1(csr_asyn_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(tstmx2_to_tstmx0), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(tstmx4_to_tstmx2), .shift_en(csr_actreden[10]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0157), .odat1_aib(net0340),
     .jtag_rx_scan_out(jtag_rx_scan_in_12x6), .odat0_aib(net0339),
     .oclk_aib(net0337), .last_bs_out(last_bs_in_12x6),
     .oclkb_aib(net0338), .jtag_clkdr_in(jtag_clkdr_in6r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_11x6),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_11x6), .iopad(iopad_tstmx[2]),
     .oclkn(net0336), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xtstmx3 ( .idata1_in1_jtag_out(net0819),
     .async_dat_in1_jtag_out(net0710), .idata0_in1_jtag_out(net0781),
     .prev_io_shift_en(csr_actreden[9]), .jtag_clkdr_outn(net0516),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(jtag_intest), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(jtag_rstb_en), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0354), .oclk_out(net0343), .oclkb_out(net0344),
     .odat0_out(net0345), .odat1_out(net0346),
     .odat_async_out(tstmx[3]), .pd_data_out(net0347),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0(csr_asyn_rxen_int[2:0]),
     .irxen_in1(csr_asyn_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(tstmx3_to_tstmx1), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(tstmx5_to_tstmx3), .shift_en(csr_actreden[10]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0152), .odat1_aib(net0352),
     .jtag_rx_scan_out(jtag_rx_scan_in_12x5), .odat0_aib(net0351),
     .oclk_aib(net0349), .last_bs_out(last_bs_in_12x5),
     .oclkb_aib(net0350), .jtag_clkdr_in(jtag_clkdr_in5r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_11x5),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_11x5), .iopad(iopad_tstmx[3]),
     .oclkn(net0348), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xio_oe0 ( .idata1_in1_jtag_out(net0785),
     .async_dat_in1_jtag_out(net0782), .idata0_in1_jtag_out(net0717),
     .prev_io_shift_en(csr_actreden[7]), .jtag_clkdr_outn(net0517),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(jtag_intest), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(jtag_rstb_en), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0366), .oclk_out(net0355), .oclkb_out(net0356),
     .odat0_out(net0357), .odat1_out(net0358),
     .odat_async_out(io_out[6]), .pd_data_out(net0359),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0(csr_asyn_rxen_int[2:0]),
     .irxen_in1(csr_asyn_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(out6_to_out4), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(tstmx0_to_out6), .shift_en(csr_actreden[8]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0618), .odat1_aib(net0364),
     .jtag_rx_scan_out(jtag_rx_scan_in_10x6), .odat0_aib(net0363),
     .oclk_aib(net0361), .last_bs_out(last_bs_in_10x6),
     .oclkb_aib(net0362), .jtag_clkdr_in(jtag_clkdr_in6r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_09x6),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_09x6), .iopad(iopad_io_out[6]),
     .oclkn(net0360), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xio_oe1 ( .idata1_in1_jtag_out(net0759),
     .async_dat_in1_jtag_out(net0813), .idata0_in1_jtag_out(net0741),
     .prev_io_shift_en(csr_actreden[7]), .jtag_clkdr_outn(net0518),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(jtag_intest), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(jtag_rstb_en), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0378), .oclk_out(net0367), .oclkb_out(net0368),
     .odat0_out(net0369), .odat1_out(net0370),
     .odat_async_out(io_out[7]), .pd_data_out(net0371),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0(csr_asyn_rxen_int[2:0]),
     .irxen_in1(csr_asyn_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(out7_to_out5), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(tstmx1_to_out7), .shift_en(csr_actreden[8]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0715), .odat1_aib(net0376),
     .jtag_rx_scan_out(jtag_rx_scan_in_10x5), .odat0_aib(net0375),
     .oclk_aib(net0373), .last_bs_out(last_bs_in_10x5),
     .oclkb_aib(net0374), .jtag_clkdr_in(jtag_clkdr_in5r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_09x5),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_09x5), .iopad(iopad_io_out[7]),
     .oclkn(net0372), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xtstmx0 ( .idata1_in1_jtag_out(net0791),
     .async_dat_in1_jtag_out(net0783), .idata0_in1_jtag_out(net0803),
     .prev_io_shift_en(csr_actreden[8]), .jtag_clkdr_outn(net0519),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(jtag_intest), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(jtag_rstb_en), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0223), .oclk_out(net0488), .oclkb_out(net0489),
     .odat0_out(net0474), .odat1_out(net0215),
     .odat_async_out(tstmx[0]), .pd_data_out(net0216),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0(csr_asyn_rxen_int[2:0]),
     .irxen_in1(csr_asyn_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(tstmx0_to_out6), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(tstmx2_to_tstmx0), .shift_en(csr_actreden[9]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0632), .odat1_aib(net0221),
     .jtag_rx_scan_out(jtag_rx_scan_in_11x6), .odat0_aib(net0220),
     .oclk_aib(net0218), .last_bs_out(last_bs_in_11x6),
     .oclkb_aib(net0219), .jtag_clkdr_in(jtag_clkdr_in6r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_10x6),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_10x6), .iopad(iopad_tstmx[0]),
     .oclkn(net0217), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xtstmx1 ( .idata1_in1_jtag_out(net0761),
     .async_dat_in1_jtag_out(net0690), .idata0_in1_jtag_out(net0794),
     .prev_io_shift_en(csr_actreden[8]), .jtag_clkdr_outn(net0520),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(jtag_intest), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(jtag_rstb_en), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0235), .oclk_out(net0224), .oclkb_out(net0225),
     .odat0_out(net0226), .odat1_out(net0227),
     .odat_async_out(tstmx[1]), .pd_data_out(net0228),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0(csr_asyn_rxen_int[2:0]),
     .irxen_in1(csr_asyn_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(tstmx1_to_out7), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(tstmx3_to_tstmx1), .shift_en(csr_actreden[9]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0721), .odat1_aib(net0233),
     .jtag_rx_scan_out(jtag_rx_scan_in_11x5), .odat0_aib(net0487),
     .oclk_aib(net0485), .last_bs_out(last_bs_in_11x5),
     .oclkb_aib(net0231), .jtag_clkdr_in(jtag_clkdr_in5r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_10x5),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_10x5), .iopad(iopad_tstmx[1]),
     .oclkn(net0229), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xtstmx6 ( .idata1_in1_jtag_out(net0636),
     .async_dat_in1_jtag_out(net0784), .idata0_in1_jtag_out(net0638),
     .prev_io_shift_en(csr_actreden[11]), .jtag_clkdr_outn(net0521),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(jtag_intest), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(jtag_rstb_en), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0247), .oclk_out(net0236), .oclkb_out(net0237),
     .odat0_out(net0238), .odat1_out(net0239),
     .odat_async_out(tstmx[6]), .pd_data_out(net0240),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0(csr_asyn_rxen_int[2:0]),
     .irxen_in1(csr_asyn_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(tstmx6_to_tstmx4), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(auxactred1_to_tstmx6),
     .shift_en(csr_actreden[12]), .pd_data_in1(vssl_aibndaux),
     .dig_rstb(dig_rstb), .jtag_clkdr_out(net0161),
     .odat1_aib(net0245), .jtag_rx_scan_out(jtag_rx_scan_in_11x8),
     .odat0_aib(net0244), .oclk_aib(net0242),
     .last_bs_out(last_bs_in_11x8), .oclkb_aib(net0243),
     .jtag_clkdr_in(jtag_clkdr_in8r), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_in_12x8),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_12x8), .iopad(iopad_tstmx[6]),
     .oclkn(net0241), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xtstmx7 ( .idata1_in1_jtag_out(net0642),
     .async_dat_in1_jtag_out(net0733), .idata0_in1_jtag_out(net0716),
     .prev_io_shift_en(csr_actreden[11]), .jtag_clkdr_outn(net0522),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(jtag_intest), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(jtag_rstb_en), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0259), .oclk_out(net0248), .oclkb_out(net0249),
     .odat0_out(net0250), .odat1_out(net0251),
     .odat_async_out(tstmx[7]), .pd_data_out(net0252),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0(csr_asyn_rxen_int[2:0]),
     .irxen_in1(csr_asyn_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(tstmx7_to_tstmx5), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(auxactred2_to_tstmx7),
     .shift_en(csr_actreden[12]), .pd_data_in1(vssl_aibndaux),
     .dig_rstb(dig_rstb), .jtag_clkdr_out(net0156),
     .odat1_aib(net0257), .jtag_rx_scan_out(jtag_rx_scan_in_11x7),
     .odat0_aib(net0256), .oclk_aib(net0254),
     .last_bs_out(last_bs_in_11x7), .oclkb_aib(net0255),
     .jtag_clkdr_in(jtag_clkdr_in7r), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_in_12x7),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_12x7), .iopad(iopad_tstmx[7]),
     .oclkn(net0253), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xio_in6 ( .idata1_in1_jtag_out(net0676),
     .async_dat_in1_jtag_out(net0724), .idata0_in1_jtag_out(net0797),
     .prev_io_shift_en(csr_actreden[6]), .jtag_clkdr_outn(net0523),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(jtag_intest), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(jtag_rstb_en), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0271), .oclk_out(net0260), .oclkb_out(net0261),
     .odat0_out(net0262), .odat1_out(net0263),
     .odat_async_out(io_out[4]), .pd_data_out(net0264),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0(csr_asyn_rxen_int[2:0]),
     .irxen_in1(csr_asyn_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(out4_to_out2), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(out6_to_out4), .shift_en(csr_actreden[7]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0695), .odat1_aib(net0269),
     .jtag_rx_scan_out(jtag_rx_scan_in_09x6), .odat0_aib(net0268),
     .oclk_aib(net0266), .last_bs_out(last_bs_in_09x6),
     .oclkb_aib(net0267), .jtag_clkdr_in(jtag_clkdr_in6r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_08x6),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_08x6), .iopad(iopad_io_out[4]),
     .oclkn(net0265), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xio_in7 ( .idata1_in1_jtag_out(net0802),
     .async_dat_in1_jtag_out(net0688), .idata0_in1_jtag_out(net0817),
     .prev_io_shift_en(csr_actreden[6]), .jtag_clkdr_outn(net0524),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(jtag_intest), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(jtag_rstb_en), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0283), .oclk_out(net0272), .oclkb_out(net0273),
     .odat0_out(net0274), .odat1_out(net0275),
     .odat_async_out(io_out[5]), .pd_data_out(net0276),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0(csr_asyn_rxen_int[2:0]),
     .irxen_in1(csr_asyn_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(out5_to_out3), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(out7_to_out5), .shift_en(csr_actreden[7]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0703), .odat1_aib(net0281),
     .jtag_rx_scan_out(jtag_rx_scan_in_09x5), .odat0_aib(net0280),
     .oclk_aib(net0278), .last_bs_out(last_bs_in_09x5),
     .oclkb_aib(net0279), .jtag_clkdr_in(jtag_clkdr_in5r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_08x5),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_08x5), .iopad(iopad_io_out[5]),
     .oclkn(net0277), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xio_in4 ( .idata1_in1_jtag_out(net0234),
     .async_dat_in1_jtag_out(net0766), .idata0_in1_jtag_out(net0809),
     .prev_io_shift_en(csr_actreden[5]), .jtag_clkdr_outn(net0525),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(jtag_intest), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(jtag_rstb_en), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0295), .oclk_out(net0284), .oclkb_out(net0285),
     .odat0_out(net0286), .odat1_out(net0287),
     .odat_async_out(io_out[2]), .pd_data_out(net0288),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0(csr_asyn_rxen_int[2:0]),
     .irxen_in1(csr_asyn_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(out2_to_out0), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(out4_to_out2), .shift_en(csr_actreden[6]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0687), .odat1_aib(net0293),
     .jtag_rx_scan_out(jtag_rx_scan_in_08x6), .odat0_aib(net0292),
     .oclk_aib(net0290), .last_bs_out(last_bs_in_08x6),
     .oclkb_aib(net0291), .jtag_clkdr_in(jtag_clkdr_in6r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_07x6),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_07x6), .iopad(iopad_io_out[2]),
     .oclkn(net0289), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xio_in5 ( .idata1_in1_jtag_out(net0763),
     .async_dat_in1_jtag_out(net0712), .idata0_in1_jtag_out(net0812),
     .prev_io_shift_en(csr_actreden[5]), .jtag_clkdr_outn(net0526),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(jtag_intest), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(jtag_rstb_en), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0469), .oclk_out(net0296), .oclkb_out(net0297),
     .odat0_out(net0298), .odat1_out(net0299),
     .odat_async_out(io_out[3]), .pd_data_out(net0479),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0(csr_asyn_rxen_int[2:0]),
     .irxen_in1(csr_asyn_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(out3_to_out1), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(out5_to_out3), .shift_en(csr_actreden[6]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0727), .odat1_aib(net0305),
     .jtag_rx_scan_out(jtag_rx_scan_in_08x5), .odat0_aib(net0480),
     .oclk_aib(net0477), .last_bs_out(last_bs_in_08x5),
     .oclkb_aib(net0303), .jtag_clkdr_in(jtag_clkdr_in5r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_07x5),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_07x5), .iopad(iopad_io_out[3]),
     .oclkn(net0481), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xio_in2 ( .idata1_in1_jtag_out(net0765),
     .async_dat_in1_jtag_out(net0821), .idata0_in1_jtag_out(net0737),
     .prev_io_shift_en(csr_actreden[4]), .jtag_clkdr_outn(net0527),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(jtag_intest), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(jtag_rstb_en), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0319), .oclk_out(net0482), .oclkb_out(net0309),
     .odat0_out(net0473), .odat1_out(net0311),
     .odat_async_out(io_out[0]), .pd_data_out(net0312),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(oe0_to_out0),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(csr_asyn_dataselb),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1(csr_asyn_ndrv_int[1:0]), .ipdrv_in0({vssl_aibndaux,
     vssl_aibndaux}), .ipdrv_in1(csr_asyn_pdrv_int[1:0]),
     .irxen_in0(csr_asyn_rxen_int[2:0]), .irxen_in1({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(csr_asyn_txen_int), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net0318), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(out2_to_out0), .shift_en(csr_actreden[5]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0613), .odat1_aib(net0472),
     .jtag_rx_scan_out(jtag_rx_scan_in_07x6), .odat0_aib(net0483),
     .oclk_aib(net0314), .last_bs_out(last_bs_in_07x6),
     .oclkb_aib(net0471), .jtag_clkdr_in(jtag_clkdr_in6l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_06x6),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_06x6), .iopad(iopad_io_out[0]),
     .oclkn(net0478), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xio_in3 ( .idata1_in1_jtag_out(net0778),
     .async_dat_in1_jtag_out(net0739), .idata0_in1_jtag_out(net0764),
     .prev_io_shift_en(csr_actreden[4]), .jtag_clkdr_outn(net0528),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(jtag_intest), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(jtag_rstb_en), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0331), .oclk_out(net0320), .oclkb_out(net0321),
     .odat0_out(net0322), .odat1_out(net0323),
     .odat_async_out(io_out[1]), .pd_data_out(net0324),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(oe1_to_out1),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(csr_asyn_dataselb),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1(csr_asyn_ndrv_int[1:0]), .ipdrv_in0({vssl_aibndaux,
     vssl_aibndaux}), .ipdrv_in1(csr_asyn_pdrv_int[1:0]),
     .irxen_in0(csr_asyn_rxen_int[2:0]), .irxen_in1({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(csr_asyn_txen_int), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net0330), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(out3_to_out1), .shift_en(csr_actreden[5]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0583), .odat1_aib(net0329),
     .jtag_rx_scan_out(jtag_rx_scan_in_07x5), .odat0_aib(net0328),
     .oclk_aib(net0326), .last_bs_out(last_bs_in_07x5),
     .oclkb_aib(net0327), .jtag_clkdr_in(jtag_clkdr_in5l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_06x5),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_06x5), .iopad(iopad_io_out[1]),
     .oclkn(net0325), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xio_in1 ( .idata1_in1_jtag_out(net0830),
     .async_dat_in1_jtag_out(oe1_to_out1),
     .idata0_in1_jtag_out(net0828), .prev_io_shift_en(csr_actreden[3]),
     .jtag_clkdr_outn(net0529), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibndaux), .jtag_intest(jtag_intest),
     .vccl_aibnd(vccl_aibndaux), .jtag_rstb_en(jtag_rstb_en),
     .anlg_rstb(anlg_rstb), .pd_data_aib(net0232), .oclk_out(net077),
     .oclkb_out(net078), .odat0_out(net079), .odat1_out(net080),
     .odat_async_out(net0143), .pd_data_out(net081),
     .async_dat_in0(io_oe[1]), .async_dat_in1(in7_to_oe1),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(csr_asyn_dataselb),
     .idataselb_in1(csr_asyn_dataselb), .iddren_in0(vssl_aibndaux),
     .iddren_in1(vssl_aibndaux), .ilaunch_clk_in0(vssl_aibndaux),
     .ilaunch_clk_in1(vssl_aibndaux), .ilpbk_dat_in0(vssl_aibndaux),
     .ilpbk_dat_in1(vssl_aibndaux), .ilpbk_en_in0(vssl_aibndaux),
     .ilpbk_en_in1(vssl_aibndaux), .indrv_in0(csr_asyn_ndrv_int[1:0]),
     .indrv_in1(csr_asyn_ndrv_int[1:0]),
     .ipdrv_in0(csr_asyn_pdrv_int[1:0]),
     .ipdrv_in1(csr_asyn_pdrv_int[1:0]), .irxen_in0({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .irxen_in1({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(csr_asyn_txen_int),
     .itxen_in1(csr_asyn_txen_int), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net087), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(csr_actreden[4]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0711), .odat1_aib(net086),
     .jtag_rx_scan_out(jtag_rx_scan_in_06x5), .odat0_aib(net085),
     .oclk_aib(net083), .last_bs_out(last_bs_in_06x5),
     .oclkb_aib(net084), .jtag_clkdr_in(jtag_clkdr_in5l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_05x5),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_05x5), .iopad(iopad_io_oe[1]),
     .oclkn(net082), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xio_in0 ( .idata1_in1_jtag_out(net0780),
     .async_dat_in1_jtag_out(oe0_to_out0),
     .idata0_in1_jtag_out(net0826), .prev_io_shift_en(csr_actreden[3]),
     .jtag_clkdr_outn(net0530), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibndaux), .jtag_intest(jtag_intest),
     .vccl_aibnd(vccl_aibndaux), .jtag_rstb_en(jtag_rstb_en),
     .anlg_rstb(anlg_rstb), .pd_data_aib(net0317), .oclk_out(net0166),
     .oclkb_out(net0167), .odat0_out(net0214), .odat1_out(net0230),
     .odat_async_out(net0144), .pd_data_out(net0169),
     .async_dat_in0(io_oe[0]), .async_dat_in1(in6_to_oe0),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(csr_asyn_dataselb),
     .idataselb_in1(csr_asyn_dataselb), .iddren_in0(vssl_aibndaux),
     .iddren_in1(vssl_aibndaux), .ilaunch_clk_in0(vssl_aibndaux),
     .ilaunch_clk_in1(vssl_aibndaux), .ilpbk_dat_in0(vssl_aibndaux),
     .ilpbk_dat_in1(vssl_aibndaux), .ilpbk_en_in0(vssl_aibndaux),
     .ilpbk_en_in1(vssl_aibndaux), .indrv_in0(csr_asyn_ndrv_int[1:0]),
     .indrv_in1(csr_asyn_ndrv_int[1:0]),
     .ipdrv_in0(csr_asyn_pdrv_int[1:0]),
     .ipdrv_in1(csr_asyn_pdrv_int[1:0]), .irxen_in0({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .irxen_in1({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(csr_asyn_txen_int),
     .itxen_in1(csr_asyn_txen_int), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net0313), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(csr_actreden[4]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0684), .odat1_aib(net0304),
     .jtag_rx_scan_out(jtag_rx_scan_in_06x6), .odat0_aib(net0300),
     .oclk_aib(net0315), .last_bs_out(last_bs_in_06x6),
     .oclkb_aib(net0310), .jtag_clkdr_in(jtag_clkdr_in6l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_05x6),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_05x6), .iopad(iopad_io_oe[0]),
     .oclkn(net0170), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xio_out6 ( .idata1_in1_jtag_out(net0679),
     .async_dat_in1_jtag_out(in6_to_oe0),
     .idata0_in1_jtag_out(net0829), .prev_io_shift_en(csr_actreden[2]),
     .jtag_clkdr_outn(net0531), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibndaux), .jtag_intest(jtag_intest),
     .vccl_aibnd(vccl_aibndaux), .jtag_rstb_en(jtag_rstb_en),
     .anlg_rstb(anlg_rstb), .pd_data_aib(net0308), .oclk_out(net0301),
     .oclkb_out(net0189), .odat0_out(net0190), .odat1_out(net0191),
     .odat_async_out(net0192), .pd_data_out(net0307),
     .async_dat_in0(io_in[6]), .async_dat_in1(in4_to_in6),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(csr_asyn_dataselb),
     .idataselb_in1(csr_asyn_dataselb), .iddren_in0(vssl_aibndaux),
     .iddren_in1(vssl_aibndaux), .ilaunch_clk_in0(vssl_aibndaux),
     .ilaunch_clk_in1(vssl_aibndaux), .ilpbk_dat_in0(vssl_aibndaux),
     .ilpbk_dat_in1(vssl_aibndaux), .ilpbk_en_in0(vssl_aibndaux),
     .ilpbk_en_in1(vssl_aibndaux), .indrv_in0(csr_asyn_ndrv_int[1:0]),
     .indrv_in1(csr_asyn_ndrv_int[1:0]),
     .ipdrv_in0(csr_asyn_pdrv_int[1:0]),
     .ipdrv_in1(csr_asyn_pdrv_int[1:0]), .irxen_in0({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .irxen_in1({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(csr_asyn_txen_int),
     .itxen_in1(csr_asyn_txen_int), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net0316), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(csr_actreden[3]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0696), .odat1_aib(net0198),
     .jtag_rx_scan_out(jtag_rx_scan_in_05x6), .odat0_aib(net0306),
     .oclk_aib(net0302), .last_bs_out(last_bs_in_05x6),
     .oclkb_aib(net0196), .jtag_clkdr_in(jtag_clkdr_in6l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_04x6),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_04x6), .iopad(iopad_io_in[6]),
     .oclkn(net0194), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xio_out7 ( .idata1_in1_jtag_out(net0155),
     .async_dat_in1_jtag_out(in7_to_oe1),
     .idata0_in1_jtag_out(net0154), .prev_io_shift_en(csr_actreden[2]),
     .jtag_clkdr_outn(net0532), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibndaux), .jtag_intest(jtag_intest),
     .vccl_aibnd(vccl_aibndaux), .jtag_rstb_en(jtag_rstb_en),
     .anlg_rstb(anlg_rstb), .pd_data_aib(net0213), .oclk_out(net0201),
     .oclkb_out(net0202), .odat0_out(net0203), .odat1_out(net0204),
     .odat_async_out(net0205), .pd_data_out(net0206),
     .async_dat_in0(io_in[7]), .async_dat_in1(in5_to_in7),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(csr_asyn_dataselb),
     .idataselb_in1(csr_asyn_dataselb), .iddren_in0(vssl_aibndaux),
     .iddren_in1(vssl_aibndaux), .ilaunch_clk_in0(vssl_aibndaux),
     .ilaunch_clk_in1(vssl_aibndaux), .ilpbk_dat_in0(vssl_aibndaux),
     .ilpbk_dat_in1(vssl_aibndaux), .ilpbk_en_in0(vssl_aibndaux),
     .ilpbk_en_in1(vssl_aibndaux), .indrv_in0(csr_asyn_ndrv_int[1:0]),
     .indrv_in1(csr_asyn_ndrv_int[1:0]),
     .ipdrv_in0(csr_asyn_pdrv_int[1:0]),
     .ipdrv_in1(csr_asyn_pdrv_int[1:0]), .irxen_in0({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .irxen_in1({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(csr_asyn_txen_int),
     .itxen_in1(csr_asyn_txen_int), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net0212), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(csr_actreden[3]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0726), .odat1_aib(net0211),
     .jtag_rx_scan_out(jtag_rx_scan_in_05x5), .odat0_aib(net0210),
     .oclk_aib(net0208), .last_bs_out(last_bs_in_05x5),
     .oclkb_aib(net0209), .jtag_clkdr_in(jtag_clkdr_in5l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_04x5),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_04x5), .iopad(iopad_io_in[7]),
     .oclkn(net0207), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xio_out4 ( .idata1_in1_jtag_out(net0816),
     .async_dat_in1_jtag_out(in4_to_in6),
     .idata0_in1_jtag_out(net0694), .prev_io_shift_en(csr_actreden[1]),
     .jtag_clkdr_outn(net0533), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibndaux), .jtag_intest(jtag_intest),
     .vccl_aibnd(vccl_aibndaux), .jtag_rstb_en(jtag_rstb_en),
     .anlg_rstb(anlg_rstb), .pd_data_aib(net0101), .oclk_out(net088),
     .oclkb_out(net089), .odat0_out(net090), .odat1_out(net091),
     .odat_async_out(net092), .pd_data_out(net093),
     .async_dat_in0(io_in[4]), .async_dat_in1(in2_to_in4),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(csr_asyn_dataselb),
     .idataselb_in1(csr_asyn_dataselb), .iddren_in0(vssl_aibndaux),
     .iddren_in1(vssl_aibndaux), .ilaunch_clk_in0(vssl_aibndaux),
     .ilaunch_clk_in1(vssl_aibndaux), .ilpbk_dat_in0(vssl_aibndaux),
     .ilpbk_dat_in1(vssl_aibndaux), .ilpbk_en_in0(vssl_aibndaux),
     .ilpbk_en_in1(vssl_aibndaux), .indrv_in0(csr_asyn_ndrv_int[1:0]),
     .indrv_in1(csr_asyn_ndrv_int[1:0]),
     .ipdrv_in0(csr_asyn_pdrv_int[1:0]),
     .ipdrv_in1(csr_asyn_pdrv_int[1:0]), .irxen_in0({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .irxen_in1({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(csr_asyn_txen_int),
     .itxen_in1(csr_asyn_txen_int), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net0100), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(csr_actreden[2]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0610), .odat1_aib(net099),
     .jtag_rx_scan_out(jtag_rx_scan_in_04x6), .odat0_aib(net098),
     .oclk_aib(net096), .last_bs_out(last_bs_in_04x6),
     .oclkb_aib(net097), .jtag_clkdr_in(jtag_clkdr_in6l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_03x6),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_03x6), .iopad(iopad_io_in[4]),
     .oclkn(net095), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xio_out5 ( .idata1_in1_jtag_out(net0648),
     .async_dat_in1_jtag_out(in5_to_in7),
     .idata0_in1_jtag_out(net0770), .prev_io_shift_en(csr_actreden[1]),
     .jtag_clkdr_outn(net0534), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibndaux), .jtag_intest(jtag_intest),
     .vccl_aibnd(vccl_aibndaux), .jtag_rstb_en(jtag_rstb_en),
     .anlg_rstb(anlg_rstb), .pd_data_aib(net0188), .oclk_out(net094),
     .oclkb_out(net0102), .odat0_out(net0195), .odat1_out(net0185),
     .odat_async_out(net0181), .pd_data_out(net0182),
     .async_dat_in0(io_in[5]), .async_dat_in1(in3_to_in5),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(csr_asyn_dataselb),
     .idataselb_in1(csr_asyn_dataselb), .iddren_in0(vssl_aibndaux),
     .iddren_in1(vssl_aibndaux), .ilaunch_clk_in0(vssl_aibndaux),
     .ilaunch_clk_in1(vssl_aibndaux), .ilpbk_dat_in0(vssl_aibndaux),
     .ilpbk_dat_in1(vssl_aibndaux), .ilpbk_en_in0(vssl_aibndaux),
     .ilpbk_en_in1(vssl_aibndaux), .indrv_in0(csr_asyn_ndrv_int[1:0]),
     .indrv_in1(csr_asyn_ndrv_int[1:0]),
     .ipdrv_in0(csr_asyn_pdrv_int[1:0]),
     .ipdrv_in1(csr_asyn_pdrv_int[1:0]), .irxen_in0({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .irxen_in1({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(csr_asyn_txen_int),
     .itxen_in1(csr_asyn_txen_int), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net0200), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(csr_actreden[2]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0168), .odat1_aib(net0197),
     .jtag_rx_scan_out(jtag_rx_scan_in_04x5), .odat0_aib(net0199),
     .oclk_aib(net0180), .last_bs_out(last_bs_in_04x5),
     .oclkb_aib(net0193), .jtag_clkdr_in(jtag_clkdr_in5l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_03x5),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_03x5), .iopad(iopad_io_in[5]),
     .oclkn(net0184), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xio_out2 ( .idata1_in1_jtag_out(net0827),
     .async_dat_in1_jtag_out(in2_to_in4),
     .idata0_in1_jtag_out(net0750), .prev_io_shift_en(csr_actreden[0]),
     .jtag_clkdr_outn(net0535), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibndaux), .jtag_intest(jtag_intest),
     .vccl_aibnd(vccl_aibndaux), .jtag_rstb_en(jtag_rstb_en),
     .anlg_rstb(anlg_rstb), .pd_data_aib(net0115), .oclk_out(net0103),
     .oclkb_out(net0104), .odat0_out(net0105), .odat1_out(net0106),
     .odat_async_out(net0107), .pd_data_out(net0108),
     .async_dat_in0(io_in[2]), .async_dat_in1(in0_to_in2),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(csr_asyn_dataselb),
     .idataselb_in1(csr_asyn_dataselb), .iddren_in0(vssl_aibndaux),
     .iddren_in1(vssl_aibndaux), .ilaunch_clk_in0(vssl_aibndaux),
     .ilaunch_clk_in1(vssl_aibndaux), .ilpbk_dat_in0(vssl_aibndaux),
     .ilpbk_dat_in1(vssl_aibndaux), .ilpbk_en_in0(vssl_aibndaux),
     .ilpbk_en_in1(vssl_aibndaux), .indrv_in0(csr_asyn_ndrv_int[1:0]),
     .indrv_in1(csr_asyn_ndrv_int[1:0]),
     .ipdrv_in0(csr_asyn_pdrv_int[1:0]),
     .ipdrv_in1(csr_asyn_pdrv_int[1:0]), .irxen_in0({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .irxen_in1({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(csr_asyn_txen_int),
     .itxen_in1(csr_asyn_txen_int), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net0114), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(csr_actreden[1]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0590), .odat1_aib(net0113),
     .jtag_rx_scan_out(jtag_rx_scan_in_03x6), .odat0_aib(net0112),
     .oclk_aib(net0110), .last_bs_out(last_bs_in_03x6),
     .oclkb_aib(net0111), .jtag_clkdr_in(jtag_clkdr_in6l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_02x6),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_02x6), .iopad(iopad_io_in[2]),
     .oclkn(net0109), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xio_out3 ( .idata1_in1_jtag_out(net0159),
     .async_dat_in1_jtag_out(in3_to_in5),
     .idata0_in1_jtag_out(net0158), .prev_io_shift_en(csr_actreden[0]),
     .jtag_clkdr_outn(net0536), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibndaux), .jtag_intest(jtag_intest),
     .vccl_aibnd(vccl_aibndaux), .jtag_rstb_en(jtag_rstb_en),
     .anlg_rstb(anlg_rstb), .pd_data_aib(net0176), .oclk_out(net0116),
     .oclkb_out(net0117), .odat0_out(net0172), .odat1_out(net0177),
     .odat_async_out(net0118), .pd_data_out(net0119),
     .async_dat_in0(io_in[3]), .async_dat_in1(in1_to_in3),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(csr_asyn_dataselb),
     .idataselb_in1(csr_asyn_dataselb), .iddren_in0(vssl_aibndaux),
     .iddren_in1(vssl_aibndaux), .ilaunch_clk_in0(vssl_aibndaux),
     .ilaunch_clk_in1(vssl_aibndaux), .ilpbk_dat_in0(vssl_aibndaux),
     .ilpbk_dat_in1(vssl_aibndaux), .ilpbk_en_in0(vssl_aibndaux),
     .ilpbk_en_in1(vssl_aibndaux), .indrv_in0(csr_asyn_ndrv_int[1:0]),
     .indrv_in1(csr_asyn_ndrv_int[1:0]),
     .ipdrv_in0(csr_asyn_pdrv_int[1:0]),
     .ipdrv_in1(csr_asyn_pdrv_int[1:0]), .irxen_in0({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .irxen_in1({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(csr_asyn_txen_int),
     .itxen_in1(csr_asyn_txen_int), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net0173), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(csr_actreden[1]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0165), .odat1_aib(net0171),
     .jtag_rx_scan_out(jtag_rx_scan_in_03x5), .odat0_aib(net0123),
     .oclk_aib(net0121), .last_bs_out(last_bs_in_03x5),
     .oclkb_aib(net0122), .jtag_clkdr_in(jtag_clkdr_in5l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_in_02x5),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_02x5), .iopad(iopad_io_in[3]),
     .oclkn(net0120), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xio_out0 ( .idata1_in1_jtag_out(net0796),
     .async_dat_in1_jtag_out(in0_to_in2),
     .idata0_in1_jtag_out(net0814), .prev_io_shift_en(vssl_aibndaux),
     .jtag_clkdr_outn(net0537), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibndaux), .jtag_intest(jtag_intest),
     .vccl_aibnd(vccl_aibndaux), .jtag_rstb_en(jtag_rstb_en),
     .anlg_rstb(anlg_rstb), .pd_data_aib(net0130), .oclk_out(net0442),
     .oclkb_out(net0416), .odat0_out(net028), .odat1_out(net029),
     .odat_async_out(net0385), .pd_data_out(net0402),
     .async_dat_in0(io_in[0]), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(csr_asyn_dataselb), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0(csr_asyn_ndrv_int[1:0]),
     .indrv_in1(csr_asyn_ndrv_int[1:0]),
     .ipdrv_in0(csr_asyn_pdrv_int[1:0]),
     .ipdrv_in1(csr_asyn_pdrv_int[1:0]), .irxen_in0({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .irxen_in1({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(csr_asyn_txen_int),
     .itxen_in1(csr_asyn_txen_int), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net0129), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(csr_actreden[0]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0666), .odat1_aib(net0128),
     .jtag_rx_scan_out(jtag_rx_scan_in_02x6), .odat0_aib(net0127),
     .oclk_aib(net0125), .last_bs_out(last_bs_in_02x6),
     .oclkb_aib(net0126), .jtag_clkdr_in(jtag_clkdr_in6l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_tx_scan_in_01x6),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_01x6), .iopad(iopad_io_in[0]),
     .oclkn(net0124), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top  xio_out1 ( .idata1_in1_jtag_out(net0825),
     .async_dat_in1_jtag_out(in1_to_in3),
     .idata0_in1_jtag_out(net0655), .prev_io_shift_en(vssl_aibndaux),
     .jtag_clkdr_outn(net0538), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibndaux), .jtag_intest(jtag_intest),
     .vccl_aibnd(vccl_aibndaux), .jtag_rstb_en(jtag_rstb_en),
     .anlg_rstb(anlg_rstb), .pd_data_aib(net051), .oclk_out(net041),
     .oclkb_out(net042), .odat0_out(net0174), .odat1_out(net0175),
     .odat_async_out(net043), .pd_data_out(net044),
     .async_dat_in0(io_in[1]), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(csr_asyn_dataselb), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0(csr_asyn_ndrv_int[1:0]),
     .indrv_in1(csr_asyn_ndrv_int[1:0]),
     .ipdrv_in0(csr_asyn_pdrv_int[1:0]),
     .ipdrv_in1(csr_asyn_pdrv_int[1:0]), .irxen_in0({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .irxen_in1({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(csr_asyn_txen_int),
     .itxen_in1(csr_asyn_txen_int), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net050), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(csr_actreden[0]),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net0164), .odat1_aib(net049),
     .jtag_rx_scan_out(jtag_rx_scan_in_02x5), .odat0_aib(net048),
     .oclk_aib(net046), .last_bs_out(last_bs_in_02x5),
     .oclkb_aib(net047), .jtag_clkdr_in(jtag_clkdr_in5l),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_tx_scan_in_01x5),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_in_01x5), .iopad(iopad_io_in[1]),
     .oclkn(net045), .iclkn(vssl_aibndaux), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
assign csr_asyn_pdrv_int[1:0] = csr_iocsr_sel ? csr_asyn_pdrv[1:0] : {vccl_aibndaux, vssl_aibndaux};
assign csr_asyn_txen_int = csr_iocsr_sel ? csr_asyn_txen : crete_detect;
assign csr_asyn_rxen_int[2:0] = csr_iocsr_sel ? csr_asyn_rxen[2:0] : vssl_aibndaux;
assign csr_asyn_ndrv_int[1:0] = csr_iocsr_sel ? csr_asyn_ndrv[1:0] : {vccl_aibndaux, vssl_aibndaux};


endmodule

