// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. All rights reserved
// *****************************************************************************
// *****************************************************************************
//  Copyright © 2016 Altera Corporation. All rights reserved. Altera products
//  are protected under numerous U.S. and foreign patents, maskwork rights,
//  copyrights and other intellectual property laws.
// *****************************************************************************
//  Module Name :  c3lib_ecc_enc_d32_c39
//  Date        :  Tue May 24 15:08:56 2016
//  Description :  ECC encoder (based on the standard Extended Hamming Code
//                 scheme). Code generated by ecc_gen.pl script (command line
//                 options used: -num_data_bits 32).
// *****************************************************************************

module c3lib_ecc_enc_d32_c39(

  input  logic[ 31 : 0 ]	i_data,
  output logic[ 38 : 0 ]	o_code

);

assign o_code[ 0 ] = o_code[ 1 ] ^ o_code[ 2 ] ^ o_code[ 3 ] ^ o_code[ 4 ] ^ o_code[ 5 ] ^ o_code[ 6 ] ^ o_code[ 7 ] ^ o_code[ 8 ] ^ o_code[ 9 ] ^ o_code[ 10 ] ^ o_code[ 11 ] ^ o_code[ 12 ] ^ o_code[ 13 ] ^ o_code[ 14 ] ^ o_code[ 15 ] ^ o_code[ 16 ] ^ o_code[ 17 ] ^ o_code[ 18 ] ^ o_code[ 19 ] ^ o_code[ 20 ] ^ o_code[ 21 ] ^ o_code[ 22 ] ^ o_code[ 23 ] ^ o_code[ 24 ] ^ o_code[ 25 ] ^ o_code[ 26 ] ^ o_code[ 27 ] ^ o_code[ 28 ] ^ o_code[ 29 ] ^ o_code[ 30 ] ^ o_code[ 31 ] ^ o_code[ 32 ] ^ o_code[ 33 ] ^ o_code[ 34 ] ^ o_code[ 35 ] ^ o_code[ 36 ] ^ o_code[ 37 ] ^ o_code[ 38 ];
assign o_code[ 1 ] = o_code[ 3 ] ^ o_code[ 5 ] ^ o_code[ 7 ] ^ o_code[ 9 ] ^ o_code[ 11 ] ^ o_code[ 13 ] ^ o_code[ 15 ] ^ o_code[ 17 ] ^ o_code[ 19 ] ^ o_code[ 21 ] ^ o_code[ 23 ] ^ o_code[ 25 ] ^ o_code[ 27 ] ^ o_code[ 29 ] ^ o_code[ 31 ] ^ o_code[ 33 ] ^ o_code[ 35 ] ^ o_code[ 37 ];
assign o_code[ 2 ] = o_code[ 3 ] ^ o_code[ 6 ] ^ o_code[ 7 ] ^ o_code[ 10 ] ^ o_code[ 11 ] ^ o_code[ 14 ] ^ o_code[ 15 ] ^ o_code[ 18 ] ^ o_code[ 19 ] ^ o_code[ 22 ] ^ o_code[ 23 ] ^ o_code[ 26 ] ^ o_code[ 27 ] ^ o_code[ 30 ] ^ o_code[ 31 ] ^ o_code[ 34 ] ^ o_code[ 35 ] ^ o_code[ 38 ];
assign o_code[ 3 ] = i_data[ 0 ];
assign o_code[ 4 ] = o_code[ 5 ] ^ o_code[ 6 ] ^ o_code[ 7 ] ^ o_code[ 12 ] ^ o_code[ 13 ] ^ o_code[ 14 ] ^ o_code[ 15 ] ^ o_code[ 20 ] ^ o_code[ 21 ] ^ o_code[ 22 ] ^ o_code[ 23 ] ^ o_code[ 28 ] ^ o_code[ 29 ] ^ o_code[ 30 ] ^ o_code[ 31 ] ^ o_code[ 36 ] ^ o_code[ 37 ] ^ o_code[ 38 ];
assign o_code[ 5 ] = i_data[ 1 ];
assign o_code[ 6 ] = i_data[ 2 ];
assign o_code[ 7 ] = i_data[ 3 ];
assign o_code[ 8 ] = o_code[ 9 ] ^ o_code[ 10 ] ^ o_code[ 11 ] ^ o_code[ 12 ] ^ o_code[ 13 ] ^ o_code[ 14 ] ^ o_code[ 15 ] ^ o_code[ 24 ] ^ o_code[ 25 ] ^ o_code[ 26 ] ^ o_code[ 27 ] ^ o_code[ 28 ] ^ o_code[ 29 ] ^ o_code[ 30 ] ^ o_code[ 31 ];
assign o_code[ 9 ] = i_data[ 4 ];
assign o_code[ 10 ] = i_data[ 5 ];
assign o_code[ 11 ] = i_data[ 6 ];
assign o_code[ 12 ] = i_data[ 7 ];
assign o_code[ 13 ] = i_data[ 8 ];
assign o_code[ 14 ] = i_data[ 9 ];
assign o_code[ 15 ] = i_data[ 10 ];
assign o_code[ 16 ] = o_code[ 17 ] ^ o_code[ 18 ] ^ o_code[ 19 ] ^ o_code[ 20 ] ^ o_code[ 21 ] ^ o_code[ 22 ] ^ o_code[ 23 ] ^ o_code[ 24 ] ^ o_code[ 25 ] ^ o_code[ 26 ] ^ o_code[ 27 ] ^ o_code[ 28 ] ^ o_code[ 29 ] ^ o_code[ 30 ] ^ o_code[ 31 ];
assign o_code[ 17 ] = i_data[ 11 ];
assign o_code[ 18 ] = i_data[ 12 ];
assign o_code[ 19 ] = i_data[ 13 ];
assign o_code[ 20 ] = i_data[ 14 ];
assign o_code[ 21 ] = i_data[ 15 ];
assign o_code[ 22 ] = i_data[ 16 ];
assign o_code[ 23 ] = i_data[ 17 ];
assign o_code[ 24 ] = i_data[ 18 ];
assign o_code[ 25 ] = i_data[ 19 ];
assign o_code[ 26 ] = i_data[ 20 ];
assign o_code[ 27 ] = i_data[ 21 ];
assign o_code[ 28 ] = i_data[ 22 ];
assign o_code[ 29 ] = i_data[ 23 ];
assign o_code[ 30 ] = i_data[ 24 ];
assign o_code[ 31 ] = i_data[ 25 ];
assign o_code[ 32 ] = o_code[ 33 ] ^ o_code[ 34 ] ^ o_code[ 35 ] ^ o_code[ 36 ] ^ o_code[ 37 ] ^ o_code[ 38 ];
assign o_code[ 33 ] = i_data[ 26 ];
assign o_code[ 34 ] = i_data[ 27 ];
assign o_code[ 35 ] = i_data[ 28 ];
assign o_code[ 36 ] = i_data[ 29 ];
assign o_code[ 37 ] = i_data[ 30 ];
assign o_code[ 38 ] = i_data[ 31 ];

endmodule

