// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. 
module aibcr3_anaio_esd (osc_extrref);

  inout osc_extrref;

endmodule

